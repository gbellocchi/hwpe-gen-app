// ----------------------------------------------------------------------------
//
// Multi-Dataflow Composer tool - Platform Composer
// Multi-Dataflow Network module 
// Date: 2022/04/29 11:36:55
//
// ----------------------------------------------------------------------------

module multi_dataflow (
	// Input(s)
	input [7 : 0] text_data,
	input text_wr,
	output text_full,
	
	// Output(s)
	input [7 : 0] key_data,
	input key_wr,
	output key_full,
	
	// Output(s)
	input [7 : 0] rc_data,
	input rc_wr,
	output rc_full,
	
	// Output(s)
	output [7 : 0] chiped_text_data,
	output chiped_text_wr,
	input chiped_text_full,
	
	// Dynamic Parameter(s)
	
	// Monitoring
	
	// Configuration ID
	
	
	// System Signal(s)		
	input clock,
	input reset
);	

// internal signals
// ----------------------------------------------------------------------------
		


// Actors Wire(s)
	
// actor add_round_key_0
wire [127 : 0] fifo_small_add_round_key_0_in_state_data;
wire fifo_small_add_round_key_0_in_state_wr;
wire fifo_small_add_round_key_0_in_state_full;
wire [127 : 0] add_round_key_0_in_state_data;
wire add_round_key_0_in_state_rd;
wire add_round_key_0_in_state_empty;
wire [127 : 0] fifo_small_add_round_key_0_round_key_data;
wire fifo_small_add_round_key_0_round_key_wr;
wire fifo_small_add_round_key_0_round_key_full;
wire [127 : 0] add_round_key_0_round_key_data;
wire add_round_key_0_round_key_rd;
wire add_round_key_0_round_key_empty;
wire [127 : 0] add_round_key_0_out_state_data;
wire add_round_key_0_out_state_wr;
wire add_round_key_0_out_state_full;
	
// actor sub_bytes_0
wire [127 : 0] fifo_small_sub_bytes_0_in_state_data;
wire fifo_small_sub_bytes_0_in_state_wr;
wire fifo_small_sub_bytes_0_in_state_full;
wire [127 : 0] sub_bytes_0_in_state_data;
wire sub_bytes_0_in_state_rd;
wire sub_bytes_0_in_state_empty;
wire [127 : 0] sub_bytes_0_out_state_data;
wire sub_bytes_0_out_state_wr;
wire sub_bytes_0_out_state_full;
	
// actor shift_rows_0
wire [127 : 0] fifo_small_shift_rows_0_in_state_data;
wire fifo_small_shift_rows_0_in_state_wr;
wire fifo_small_shift_rows_0_in_state_full;
wire [127 : 0] shift_rows_0_in_state_data;
wire shift_rows_0_in_state_rd;
wire shift_rows_0_in_state_empty;
wire [127 : 0] shift_rows_0_out_state_data;
wire shift_rows_0_out_state_wr;
wire shift_rows_0_out_state_full;
	
// actor add_round_key_1
wire [127 : 0] fifo_small_add_round_key_1_in_state_data;
wire fifo_small_add_round_key_1_in_state_wr;
wire fifo_small_add_round_key_1_in_state_full;
wire [127 : 0] add_round_key_1_in_state_data;
wire add_round_key_1_in_state_rd;
wire add_round_key_1_in_state_empty;
wire [127 : 0] fifo_small_add_round_key_1_round_key_data;
wire fifo_small_add_round_key_1_round_key_wr;
wire fifo_small_add_round_key_1_round_key_full;
wire [127 : 0] add_round_key_1_round_key_data;
wire add_round_key_1_round_key_rd;
wire add_round_key_1_round_key_empty;
wire [127 : 0] add_round_key_1_out_state_data;
wire add_round_key_1_out_state_wr;
wire add_round_key_1_out_state_full;
	
// actor read8x16_0
wire [7 : 0] fifo_small_read8x16_0_in_token_data;
wire fifo_small_read8x16_0_in_token_wr;
wire fifo_small_read8x16_0_in_token_full;
wire [7 : 0] read8x16_0_in_token_data;
wire read8x16_0_in_token_rd;
wire read8x16_0_in_token_empty;
wire [127 : 0] read8x16_0_out_token_data;
wire read8x16_0_out_token_wr;
wire read8x16_0_out_token_full;
	
// actor read8x16_1
wire [7 : 0] fifo_small_read8x16_1_in_token_data;
wire fifo_small_read8x16_1_in_token_wr;
wire fifo_small_read8x16_1_in_token_full;
wire [7 : 0] read8x16_1_in_token_data;
wire read8x16_1_in_token_rd;
wire read8x16_1_in_token_empty;
wire [127 : 0] read8x16_1_out_token_data;
wire read8x16_1_out_token_wr;
wire read8x16_1_out_token_full;
	
// actor write16x8_0
wire [127 : 0] fifo_small_write16x8_0_in_token_data;
wire fifo_small_write16x8_0_in_token_wr;
wire fifo_small_write16x8_0_in_token_full;
wire [127 : 0] write16x8_0_in_token_data;
wire write16x8_0_in_token_rd;
wire write16x8_0_in_token_empty;
wire [7 : 0] write16x8_0_out_token_data;
wire write16x8_0_out_token_wr;
wire write16x8_0_out_token_full;
	
// actor sub_bytes_1
wire [127 : 0] fifo_small_sub_bytes_1_in_state_data;
wire fifo_small_sub_bytes_1_in_state_wr;
wire fifo_small_sub_bytes_1_in_state_full;
wire [127 : 0] sub_bytes_1_in_state_data;
wire sub_bytes_1_in_state_rd;
wire sub_bytes_1_in_state_empty;
wire [127 : 0] sub_bytes_1_out_state_data;
wire sub_bytes_1_out_state_wr;
wire sub_bytes_1_out_state_full;
	
// actor shift_rows_1
wire [127 : 0] fifo_small_shift_rows_1_in_state_data;
wire fifo_small_shift_rows_1_in_state_wr;
wire fifo_small_shift_rows_1_in_state_full;
wire [127 : 0] shift_rows_1_in_state_data;
wire shift_rows_1_in_state_rd;
wire shift_rows_1_in_state_empty;
wire [127 : 0] shift_rows_1_out_state_data;
wire shift_rows_1_out_state_wr;
wire shift_rows_1_out_state_full;
	
// actor mix_cols_0
wire [127 : 0] fifo_small_mix_cols_0_in_state_data;
wire fifo_small_mix_cols_0_in_state_wr;
wire fifo_small_mix_cols_0_in_state_full;
wire [127 : 0] mix_cols_0_in_state_data;
wire mix_cols_0_in_state_rd;
wire mix_cols_0_in_state_empty;
wire [127 : 0] mix_cols_0_out_state_data;
wire mix_cols_0_out_state_wr;
wire mix_cols_0_out_state_full;
	
// actor add_round_key_2
wire [127 : 0] fifo_small_add_round_key_2_in_state_data;
wire fifo_small_add_round_key_2_in_state_wr;
wire fifo_small_add_round_key_2_in_state_full;
wire [127 : 0] add_round_key_2_in_state_data;
wire add_round_key_2_in_state_rd;
wire add_round_key_2_in_state_empty;
wire [127 : 0] fifo_small_add_round_key_2_round_key_data;
wire fifo_small_add_round_key_2_round_key_wr;
wire fifo_small_add_round_key_2_round_key_full;
wire [127 : 0] add_round_key_2_round_key_data;
wire add_round_key_2_round_key_rd;
wire add_round_key_2_round_key_empty;
wire [127 : 0] add_round_key_2_out_state_data;
wire add_round_key_2_out_state_wr;
wire add_round_key_2_out_state_full;
	
// actor sub_bytes_2
wire [127 : 0] fifo_small_sub_bytes_2_in_state_data;
wire fifo_small_sub_bytes_2_in_state_wr;
wire fifo_small_sub_bytes_2_in_state_full;
wire [127 : 0] sub_bytes_2_in_state_data;
wire sub_bytes_2_in_state_rd;
wire sub_bytes_2_in_state_empty;
wire [127 : 0] sub_bytes_2_out_state_data;
wire sub_bytes_2_out_state_wr;
wire sub_bytes_2_out_state_full;
	
// actor shift_rows_2
wire [127 : 0] fifo_small_shift_rows_2_in_state_data;
wire fifo_small_shift_rows_2_in_state_wr;
wire fifo_small_shift_rows_2_in_state_full;
wire [127 : 0] shift_rows_2_in_state_data;
wire shift_rows_2_in_state_rd;
wire shift_rows_2_in_state_empty;
wire [127 : 0] shift_rows_2_out_state_data;
wire shift_rows_2_out_state_wr;
wire shift_rows_2_out_state_full;
	
// actor mix_cols_1
wire [127 : 0] fifo_small_mix_cols_1_in_state_data;
wire fifo_small_mix_cols_1_in_state_wr;
wire fifo_small_mix_cols_1_in_state_full;
wire [127 : 0] mix_cols_1_in_state_data;
wire mix_cols_1_in_state_rd;
wire mix_cols_1_in_state_empty;
wire [127 : 0] mix_cols_1_out_state_data;
wire mix_cols_1_out_state_wr;
wire mix_cols_1_out_state_full;
	
// actor add_round_key_3
wire [127 : 0] fifo_small_add_round_key_3_in_state_data;
wire fifo_small_add_round_key_3_in_state_wr;
wire fifo_small_add_round_key_3_in_state_full;
wire [127 : 0] add_round_key_3_in_state_data;
wire add_round_key_3_in_state_rd;
wire add_round_key_3_in_state_empty;
wire [127 : 0] fifo_small_add_round_key_3_round_key_data;
wire fifo_small_add_round_key_3_round_key_wr;
wire fifo_small_add_round_key_3_round_key_full;
wire [127 : 0] add_round_key_3_round_key_data;
wire add_round_key_3_round_key_rd;
wire add_round_key_3_round_key_empty;
wire [127 : 0] add_round_key_3_out_state_data;
wire add_round_key_3_out_state_wr;
wire add_round_key_3_out_state_full;
	
// actor sub_bytes_3
wire [127 : 0] fifo_small_sub_bytes_3_in_state_data;
wire fifo_small_sub_bytes_3_in_state_wr;
wire fifo_small_sub_bytes_3_in_state_full;
wire [127 : 0] sub_bytes_3_in_state_data;
wire sub_bytes_3_in_state_rd;
wire sub_bytes_3_in_state_empty;
wire [127 : 0] sub_bytes_3_out_state_data;
wire sub_bytes_3_out_state_wr;
wire sub_bytes_3_out_state_full;
	
// actor shift_rows_3
wire [127 : 0] fifo_small_shift_rows_3_in_state_data;
wire fifo_small_shift_rows_3_in_state_wr;
wire fifo_small_shift_rows_3_in_state_full;
wire [127 : 0] shift_rows_3_in_state_data;
wire shift_rows_3_in_state_rd;
wire shift_rows_3_in_state_empty;
wire [127 : 0] shift_rows_3_out_state_data;
wire shift_rows_3_out_state_wr;
wire shift_rows_3_out_state_full;
	
// actor mix_cols_2
wire [127 : 0] fifo_small_mix_cols_2_in_state_data;
wire fifo_small_mix_cols_2_in_state_wr;
wire fifo_small_mix_cols_2_in_state_full;
wire [127 : 0] mix_cols_2_in_state_data;
wire mix_cols_2_in_state_rd;
wire mix_cols_2_in_state_empty;
wire [127 : 0] mix_cols_2_out_state_data;
wire mix_cols_2_out_state_wr;
wire mix_cols_2_out_state_full;
	
// actor add_round_key_4
wire [127 : 0] fifo_small_add_round_key_4_in_state_data;
wire fifo_small_add_round_key_4_in_state_wr;
wire fifo_small_add_round_key_4_in_state_full;
wire [127 : 0] add_round_key_4_in_state_data;
wire add_round_key_4_in_state_rd;
wire add_round_key_4_in_state_empty;
wire [127 : 0] fifo_small_add_round_key_4_round_key_data;
wire fifo_small_add_round_key_4_round_key_wr;
wire fifo_small_add_round_key_4_round_key_full;
wire [127 : 0] add_round_key_4_round_key_data;
wire add_round_key_4_round_key_rd;
wire add_round_key_4_round_key_empty;
wire [127 : 0] add_round_key_4_out_state_data;
wire add_round_key_4_out_state_wr;
wire add_round_key_4_out_state_full;
	
// actor sub_bytes_4
wire [127 : 0] fifo_small_sub_bytes_4_in_state_data;
wire fifo_small_sub_bytes_4_in_state_wr;
wire fifo_small_sub_bytes_4_in_state_full;
wire [127 : 0] sub_bytes_4_in_state_data;
wire sub_bytes_4_in_state_rd;
wire sub_bytes_4_in_state_empty;
wire [127 : 0] sub_bytes_4_out_state_data;
wire sub_bytes_4_out_state_wr;
wire sub_bytes_4_out_state_full;
	
// actor shift_rows_4
wire [127 : 0] fifo_small_shift_rows_4_in_state_data;
wire fifo_small_shift_rows_4_in_state_wr;
wire fifo_small_shift_rows_4_in_state_full;
wire [127 : 0] shift_rows_4_in_state_data;
wire shift_rows_4_in_state_rd;
wire shift_rows_4_in_state_empty;
wire [127 : 0] shift_rows_4_out_state_data;
wire shift_rows_4_out_state_wr;
wire shift_rows_4_out_state_full;
	
// actor mix_cols_3
wire [127 : 0] fifo_small_mix_cols_3_in_state_data;
wire fifo_small_mix_cols_3_in_state_wr;
wire fifo_small_mix_cols_3_in_state_full;
wire [127 : 0] mix_cols_3_in_state_data;
wire mix_cols_3_in_state_rd;
wire mix_cols_3_in_state_empty;
wire [127 : 0] mix_cols_3_out_state_data;
wire mix_cols_3_out_state_wr;
wire mix_cols_3_out_state_full;
	
// actor add_round_key_5
wire [127 : 0] fifo_small_add_round_key_5_in_state_data;
wire fifo_small_add_round_key_5_in_state_wr;
wire fifo_small_add_round_key_5_in_state_full;
wire [127 : 0] add_round_key_5_in_state_data;
wire add_round_key_5_in_state_rd;
wire add_round_key_5_in_state_empty;
wire [127 : 0] fifo_small_add_round_key_5_round_key_data;
wire fifo_small_add_round_key_5_round_key_wr;
wire fifo_small_add_round_key_5_round_key_full;
wire [127 : 0] add_round_key_5_round_key_data;
wire add_round_key_5_round_key_rd;
wire add_round_key_5_round_key_empty;
wire [127 : 0] add_round_key_5_out_state_data;
wire add_round_key_5_out_state_wr;
wire add_round_key_5_out_state_full;
	
// actor sub_bytes_5
wire [127 : 0] fifo_small_sub_bytes_5_in_state_data;
wire fifo_small_sub_bytes_5_in_state_wr;
wire fifo_small_sub_bytes_5_in_state_full;
wire [127 : 0] sub_bytes_5_in_state_data;
wire sub_bytes_5_in_state_rd;
wire sub_bytes_5_in_state_empty;
wire [127 : 0] sub_bytes_5_out_state_data;
wire sub_bytes_5_out_state_wr;
wire sub_bytes_5_out_state_full;
	
// actor shift_rows_5
wire [127 : 0] fifo_small_shift_rows_5_in_state_data;
wire fifo_small_shift_rows_5_in_state_wr;
wire fifo_small_shift_rows_5_in_state_full;
wire [127 : 0] shift_rows_5_in_state_data;
wire shift_rows_5_in_state_rd;
wire shift_rows_5_in_state_empty;
wire [127 : 0] shift_rows_5_out_state_data;
wire shift_rows_5_out_state_wr;
wire shift_rows_5_out_state_full;
	
// actor mix_cols_4
wire [127 : 0] fifo_small_mix_cols_4_in_state_data;
wire fifo_small_mix_cols_4_in_state_wr;
wire fifo_small_mix_cols_4_in_state_full;
wire [127 : 0] mix_cols_4_in_state_data;
wire mix_cols_4_in_state_rd;
wire mix_cols_4_in_state_empty;
wire [127 : 0] mix_cols_4_out_state_data;
wire mix_cols_4_out_state_wr;
wire mix_cols_4_out_state_full;
	
// actor add_round_key_6
wire [127 : 0] fifo_small_add_round_key_6_in_state_data;
wire fifo_small_add_round_key_6_in_state_wr;
wire fifo_small_add_round_key_6_in_state_full;
wire [127 : 0] add_round_key_6_in_state_data;
wire add_round_key_6_in_state_rd;
wire add_round_key_6_in_state_empty;
wire [127 : 0] fifo_small_add_round_key_6_round_key_data;
wire fifo_small_add_round_key_6_round_key_wr;
wire fifo_small_add_round_key_6_round_key_full;
wire [127 : 0] add_round_key_6_round_key_data;
wire add_round_key_6_round_key_rd;
wire add_round_key_6_round_key_empty;
wire [127 : 0] add_round_key_6_out_state_data;
wire add_round_key_6_out_state_wr;
wire add_round_key_6_out_state_full;
	
// actor sub_bytes_6
wire [127 : 0] fifo_small_sub_bytes_6_in_state_data;
wire fifo_small_sub_bytes_6_in_state_wr;
wire fifo_small_sub_bytes_6_in_state_full;
wire [127 : 0] sub_bytes_6_in_state_data;
wire sub_bytes_6_in_state_rd;
wire sub_bytes_6_in_state_empty;
wire [127 : 0] sub_bytes_6_out_state_data;
wire sub_bytes_6_out_state_wr;
wire sub_bytes_6_out_state_full;
	
// actor shift_rows_6
wire [127 : 0] fifo_small_shift_rows_6_in_state_data;
wire fifo_small_shift_rows_6_in_state_wr;
wire fifo_small_shift_rows_6_in_state_full;
wire [127 : 0] shift_rows_6_in_state_data;
wire shift_rows_6_in_state_rd;
wire shift_rows_6_in_state_empty;
wire [127 : 0] shift_rows_6_out_state_data;
wire shift_rows_6_out_state_wr;
wire shift_rows_6_out_state_full;
	
// actor mix_cols_5
wire [127 : 0] fifo_small_mix_cols_5_in_state_data;
wire fifo_small_mix_cols_5_in_state_wr;
wire fifo_small_mix_cols_5_in_state_full;
wire [127 : 0] mix_cols_5_in_state_data;
wire mix_cols_5_in_state_rd;
wire mix_cols_5_in_state_empty;
wire [127 : 0] mix_cols_5_out_state_data;
wire mix_cols_5_out_state_wr;
wire mix_cols_5_out_state_full;
	
// actor add_round_key_7
wire [127 : 0] fifo_small_add_round_key_7_in_state_data;
wire fifo_small_add_round_key_7_in_state_wr;
wire fifo_small_add_round_key_7_in_state_full;
wire [127 : 0] add_round_key_7_in_state_data;
wire add_round_key_7_in_state_rd;
wire add_round_key_7_in_state_empty;
wire [127 : 0] fifo_small_add_round_key_7_round_key_data;
wire fifo_small_add_round_key_7_round_key_wr;
wire fifo_small_add_round_key_7_round_key_full;
wire [127 : 0] add_round_key_7_round_key_data;
wire add_round_key_7_round_key_rd;
wire add_round_key_7_round_key_empty;
wire [127 : 0] add_round_key_7_out_state_data;
wire add_round_key_7_out_state_wr;
wire add_round_key_7_out_state_full;
	
// actor sub_bytes_7
wire [127 : 0] fifo_small_sub_bytes_7_in_state_data;
wire fifo_small_sub_bytes_7_in_state_wr;
wire fifo_small_sub_bytes_7_in_state_full;
wire [127 : 0] sub_bytes_7_in_state_data;
wire sub_bytes_7_in_state_rd;
wire sub_bytes_7_in_state_empty;
wire [127 : 0] sub_bytes_7_out_state_data;
wire sub_bytes_7_out_state_wr;
wire sub_bytes_7_out_state_full;
	
// actor shift_rows_7
wire [127 : 0] fifo_small_shift_rows_7_in_state_data;
wire fifo_small_shift_rows_7_in_state_wr;
wire fifo_small_shift_rows_7_in_state_full;
wire [127 : 0] shift_rows_7_in_state_data;
wire shift_rows_7_in_state_rd;
wire shift_rows_7_in_state_empty;
wire [127 : 0] shift_rows_7_out_state_data;
wire shift_rows_7_out_state_wr;
wire shift_rows_7_out_state_full;
	
// actor mix_cols_6
wire [127 : 0] fifo_small_mix_cols_6_in_state_data;
wire fifo_small_mix_cols_6_in_state_wr;
wire fifo_small_mix_cols_6_in_state_full;
wire [127 : 0] mix_cols_6_in_state_data;
wire mix_cols_6_in_state_rd;
wire mix_cols_6_in_state_empty;
wire [127 : 0] mix_cols_6_out_state_data;
wire mix_cols_6_out_state_wr;
wire mix_cols_6_out_state_full;
	
// actor add_round_key_8
wire [127 : 0] fifo_small_add_round_key_8_in_state_data;
wire fifo_small_add_round_key_8_in_state_wr;
wire fifo_small_add_round_key_8_in_state_full;
wire [127 : 0] add_round_key_8_in_state_data;
wire add_round_key_8_in_state_rd;
wire add_round_key_8_in_state_empty;
wire [127 : 0] fifo_small_add_round_key_8_round_key_data;
wire fifo_small_add_round_key_8_round_key_wr;
wire fifo_small_add_round_key_8_round_key_full;
wire [127 : 0] add_round_key_8_round_key_data;
wire add_round_key_8_round_key_rd;
wire add_round_key_8_round_key_empty;
wire [127 : 0] add_round_key_8_out_state_data;
wire add_round_key_8_out_state_wr;
wire add_round_key_8_out_state_full;
	
// actor sub_bytes_8
wire [127 : 0] fifo_small_sub_bytes_8_in_state_data;
wire fifo_small_sub_bytes_8_in_state_wr;
wire fifo_small_sub_bytes_8_in_state_full;
wire [127 : 0] sub_bytes_8_in_state_data;
wire sub_bytes_8_in_state_rd;
wire sub_bytes_8_in_state_empty;
wire [127 : 0] sub_bytes_8_out_state_data;
wire sub_bytes_8_out_state_wr;
wire sub_bytes_8_out_state_full;
	
// actor shift_rows_8
wire [127 : 0] fifo_small_shift_rows_8_in_state_data;
wire fifo_small_shift_rows_8_in_state_wr;
wire fifo_small_shift_rows_8_in_state_full;
wire [127 : 0] shift_rows_8_in_state_data;
wire shift_rows_8_in_state_rd;
wire shift_rows_8_in_state_empty;
wire [127 : 0] shift_rows_8_out_state_data;
wire shift_rows_8_out_state_wr;
wire shift_rows_8_out_state_full;
	
// actor mix_cols_7
wire [127 : 0] fifo_small_mix_cols_7_in_state_data;
wire fifo_small_mix_cols_7_in_state_wr;
wire fifo_small_mix_cols_7_in_state_full;
wire [127 : 0] mix_cols_7_in_state_data;
wire mix_cols_7_in_state_rd;
wire mix_cols_7_in_state_empty;
wire [127 : 0] mix_cols_7_out_state_data;
wire mix_cols_7_out_state_wr;
wire mix_cols_7_out_state_full;
	
// actor add_round_key_9
wire [127 : 0] fifo_small_add_round_key_9_in_state_data;
wire fifo_small_add_round_key_9_in_state_wr;
wire fifo_small_add_round_key_9_in_state_full;
wire [127 : 0] add_round_key_9_in_state_data;
wire add_round_key_9_in_state_rd;
wire add_round_key_9_in_state_empty;
wire [127 : 0] fifo_small_add_round_key_9_round_key_data;
wire fifo_small_add_round_key_9_round_key_wr;
wire fifo_small_add_round_key_9_round_key_full;
wire [127 : 0] add_round_key_9_round_key_data;
wire add_round_key_9_round_key_rd;
wire add_round_key_9_round_key_empty;
wire [127 : 0] add_round_key_9_out_state_data;
wire add_round_key_9_out_state_wr;
wire add_round_key_9_out_state_full;
	
// actor expand_key0_128_0
wire [127 : 0] fifo_small_expand_key0_128_0_in_key_data;
wire fifo_small_expand_key0_128_0_in_key_wr;
wire fifo_small_expand_key0_128_0_in_key_full;
wire [127 : 0] expand_key0_128_0_in_key_data;
wire expand_key0_128_0_in_key_rd;
wire expand_key0_128_0_in_key_empty;
wire [7 : 0] fifo_small_expand_key0_128_0_in_rc_data;
wire fifo_small_expand_key0_128_0_in_rc_wr;
wire fifo_small_expand_key0_128_0_in_rc_full;
wire [7 : 0] expand_key0_128_0_in_rc_data;
wire expand_key0_128_0_in_rc_rd;
wire expand_key0_128_0_in_rc_empty;
wire [127 : 0] expand_key0_128_0_out_key_data;
wire expand_key0_128_0_out_key_wr;
wire expand_key0_128_0_out_key_full;
	
// actor expand_key1_128_0
wire [127 : 0] fifo_small_expand_key1_128_0_in_key_data;
wire fifo_small_expand_key1_128_0_in_key_wr;
wire fifo_small_expand_key1_128_0_in_key_full;
wire [127 : 0] expand_key1_128_0_in_key_data;
wire expand_key1_128_0_in_key_rd;
wire expand_key1_128_0_in_key_empty;
wire [127 : 0] expand_key1_128_0_out_key_data;
wire expand_key1_128_0_out_key_wr;
wire expand_key1_128_0_out_key_full;
	
// actor expand_key2_128_0
wire [127 : 0] fifo_small_expand_key2_128_0_in_key_data;
wire fifo_small_expand_key2_128_0_in_key_wr;
wire fifo_small_expand_key2_128_0_in_key_full;
wire [127 : 0] expand_key2_128_0_in_key_data;
wire expand_key2_128_0_in_key_rd;
wire expand_key2_128_0_in_key_empty;
wire [127 : 0] expand_key2_128_0_out_key_data;
wire expand_key2_128_0_out_key_wr;
wire expand_key2_128_0_out_key_full;
	
// actor expand_key3_128_0
wire [127 : 0] fifo_small_expand_key3_128_0_in_key_data;
wire fifo_small_expand_key3_128_0_in_key_wr;
wire fifo_small_expand_key3_128_0_in_key_full;
wire [127 : 0] expand_key3_128_0_in_key_data;
wire expand_key3_128_0_in_key_rd;
wire expand_key3_128_0_in_key_empty;
wire [127 : 0] expand_key3_128_0_out_key_data;
wire expand_key3_128_0_out_key_wr;
wire expand_key3_128_0_out_key_full;
	
// actor expand_key0_128_1
wire [127 : 0] fifo_small_expand_key0_128_1_in_key_data;
wire fifo_small_expand_key0_128_1_in_key_wr;
wire fifo_small_expand_key0_128_1_in_key_full;
wire [127 : 0] expand_key0_128_1_in_key_data;
wire expand_key0_128_1_in_key_rd;
wire expand_key0_128_1_in_key_empty;
wire [7 : 0] fifo_small_expand_key0_128_1_in_rc_data;
wire fifo_small_expand_key0_128_1_in_rc_wr;
wire fifo_small_expand_key0_128_1_in_rc_full;
wire [7 : 0] expand_key0_128_1_in_rc_data;
wire expand_key0_128_1_in_rc_rd;
wire expand_key0_128_1_in_rc_empty;
wire [127 : 0] expand_key0_128_1_out_key_data;
wire expand_key0_128_1_out_key_wr;
wire expand_key0_128_1_out_key_full;
	
// actor expand_key1_128_1
wire [127 : 0] fifo_small_expand_key1_128_1_in_key_data;
wire fifo_small_expand_key1_128_1_in_key_wr;
wire fifo_small_expand_key1_128_1_in_key_full;
wire [127 : 0] expand_key1_128_1_in_key_data;
wire expand_key1_128_1_in_key_rd;
wire expand_key1_128_1_in_key_empty;
wire [127 : 0] expand_key1_128_1_out_key_data;
wire expand_key1_128_1_out_key_wr;
wire expand_key1_128_1_out_key_full;
	
// actor expand_key2_128_1
wire [127 : 0] fifo_small_expand_key2_128_1_in_key_data;
wire fifo_small_expand_key2_128_1_in_key_wr;
wire fifo_small_expand_key2_128_1_in_key_full;
wire [127 : 0] expand_key2_128_1_in_key_data;
wire expand_key2_128_1_in_key_rd;
wire expand_key2_128_1_in_key_empty;
wire [127 : 0] expand_key2_128_1_out_key_data;
wire expand_key2_128_1_out_key_wr;
wire expand_key2_128_1_out_key_full;
	
// actor expand_key3_128_1
wire [127 : 0] fifo_small_expand_key3_128_1_in_key_data;
wire fifo_small_expand_key3_128_1_in_key_wr;
wire fifo_small_expand_key3_128_1_in_key_full;
wire [127 : 0] expand_key3_128_1_in_key_data;
wire expand_key3_128_1_in_key_rd;
wire expand_key3_128_1_in_key_empty;
wire [127 : 0] expand_key3_128_1_out_key_data;
wire expand_key3_128_1_out_key_wr;
wire expand_key3_128_1_out_key_full;
	
// actor expand_key0_128_2
wire [127 : 0] fifo_small_expand_key0_128_2_in_key_data;
wire fifo_small_expand_key0_128_2_in_key_wr;
wire fifo_small_expand_key0_128_2_in_key_full;
wire [127 : 0] expand_key0_128_2_in_key_data;
wire expand_key0_128_2_in_key_rd;
wire expand_key0_128_2_in_key_empty;
wire [7 : 0] fifo_small_expand_key0_128_2_in_rc_data;
wire fifo_small_expand_key0_128_2_in_rc_wr;
wire fifo_small_expand_key0_128_2_in_rc_full;
wire [7 : 0] expand_key0_128_2_in_rc_data;
wire expand_key0_128_2_in_rc_rd;
wire expand_key0_128_2_in_rc_empty;
wire [127 : 0] expand_key0_128_2_out_key_data;
wire expand_key0_128_2_out_key_wr;
wire expand_key0_128_2_out_key_full;
	
// actor expand_key1_128_2
wire [127 : 0] fifo_small_expand_key1_128_2_in_key_data;
wire fifo_small_expand_key1_128_2_in_key_wr;
wire fifo_small_expand_key1_128_2_in_key_full;
wire [127 : 0] expand_key1_128_2_in_key_data;
wire expand_key1_128_2_in_key_rd;
wire expand_key1_128_2_in_key_empty;
wire [127 : 0] expand_key1_128_2_out_key_data;
wire expand_key1_128_2_out_key_wr;
wire expand_key1_128_2_out_key_full;
	
// actor expand_key2_128_2
wire [127 : 0] fifo_small_expand_key2_128_2_in_key_data;
wire fifo_small_expand_key2_128_2_in_key_wr;
wire fifo_small_expand_key2_128_2_in_key_full;
wire [127 : 0] expand_key2_128_2_in_key_data;
wire expand_key2_128_2_in_key_rd;
wire expand_key2_128_2_in_key_empty;
wire [127 : 0] expand_key2_128_2_out_key_data;
wire expand_key2_128_2_out_key_wr;
wire expand_key2_128_2_out_key_full;
	
// actor expand_key3_128_2
wire [127 : 0] fifo_small_expand_key3_128_2_in_key_data;
wire fifo_small_expand_key3_128_2_in_key_wr;
wire fifo_small_expand_key3_128_2_in_key_full;
wire [127 : 0] expand_key3_128_2_in_key_data;
wire expand_key3_128_2_in_key_rd;
wire expand_key3_128_2_in_key_empty;
wire [127 : 0] expand_key3_128_2_out_key_data;
wire expand_key3_128_2_out_key_wr;
wire expand_key3_128_2_out_key_full;
	
// actor expand_key0_128_3
wire [127 : 0] fifo_small_expand_key0_128_3_in_key_data;
wire fifo_small_expand_key0_128_3_in_key_wr;
wire fifo_small_expand_key0_128_3_in_key_full;
wire [127 : 0] expand_key0_128_3_in_key_data;
wire expand_key0_128_3_in_key_rd;
wire expand_key0_128_3_in_key_empty;
wire [7 : 0] fifo_small_expand_key0_128_3_in_rc_data;
wire fifo_small_expand_key0_128_3_in_rc_wr;
wire fifo_small_expand_key0_128_3_in_rc_full;
wire [7 : 0] expand_key0_128_3_in_rc_data;
wire expand_key0_128_3_in_rc_rd;
wire expand_key0_128_3_in_rc_empty;
wire [127 : 0] expand_key0_128_3_out_key_data;
wire expand_key0_128_3_out_key_wr;
wire expand_key0_128_3_out_key_full;
	
// actor expand_key1_128_3
wire [127 : 0] fifo_small_expand_key1_128_3_in_key_data;
wire fifo_small_expand_key1_128_3_in_key_wr;
wire fifo_small_expand_key1_128_3_in_key_full;
wire [127 : 0] expand_key1_128_3_in_key_data;
wire expand_key1_128_3_in_key_rd;
wire expand_key1_128_3_in_key_empty;
wire [127 : 0] expand_key1_128_3_out_key_data;
wire expand_key1_128_3_out_key_wr;
wire expand_key1_128_3_out_key_full;
	
// actor expand_key2_128_3
wire [127 : 0] fifo_small_expand_key2_128_3_in_key_data;
wire fifo_small_expand_key2_128_3_in_key_wr;
wire fifo_small_expand_key2_128_3_in_key_full;
wire [127 : 0] expand_key2_128_3_in_key_data;
wire expand_key2_128_3_in_key_rd;
wire expand_key2_128_3_in_key_empty;
wire [127 : 0] expand_key2_128_3_out_key_data;
wire expand_key2_128_3_out_key_wr;
wire expand_key2_128_3_out_key_full;
	
// actor expand_key3_128_3
wire [127 : 0] fifo_small_expand_key3_128_3_in_key_data;
wire fifo_small_expand_key3_128_3_in_key_wr;
wire fifo_small_expand_key3_128_3_in_key_full;
wire [127 : 0] expand_key3_128_3_in_key_data;
wire expand_key3_128_3_in_key_rd;
wire expand_key3_128_3_in_key_empty;
wire [127 : 0] expand_key3_128_3_out_key_data;
wire expand_key3_128_3_out_key_wr;
wire expand_key3_128_3_out_key_full;
	
// actor expand_key0_128_4
wire [127 : 0] fifo_small_expand_key0_128_4_in_key_data;
wire fifo_small_expand_key0_128_4_in_key_wr;
wire fifo_small_expand_key0_128_4_in_key_full;
wire [127 : 0] expand_key0_128_4_in_key_data;
wire expand_key0_128_4_in_key_rd;
wire expand_key0_128_4_in_key_empty;
wire [7 : 0] fifo_small_expand_key0_128_4_in_rc_data;
wire fifo_small_expand_key0_128_4_in_rc_wr;
wire fifo_small_expand_key0_128_4_in_rc_full;
wire [7 : 0] expand_key0_128_4_in_rc_data;
wire expand_key0_128_4_in_rc_rd;
wire expand_key0_128_4_in_rc_empty;
wire [127 : 0] expand_key0_128_4_out_key_data;
wire expand_key0_128_4_out_key_wr;
wire expand_key0_128_4_out_key_full;
	
// actor expand_key1_128_4
wire [127 : 0] fifo_small_expand_key1_128_4_in_key_data;
wire fifo_small_expand_key1_128_4_in_key_wr;
wire fifo_small_expand_key1_128_4_in_key_full;
wire [127 : 0] expand_key1_128_4_in_key_data;
wire expand_key1_128_4_in_key_rd;
wire expand_key1_128_4_in_key_empty;
wire [127 : 0] expand_key1_128_4_out_key_data;
wire expand_key1_128_4_out_key_wr;
wire expand_key1_128_4_out_key_full;
	
// actor expand_key2_128_4
wire [127 : 0] fifo_small_expand_key2_128_4_in_key_data;
wire fifo_small_expand_key2_128_4_in_key_wr;
wire fifo_small_expand_key2_128_4_in_key_full;
wire [127 : 0] expand_key2_128_4_in_key_data;
wire expand_key2_128_4_in_key_rd;
wire expand_key2_128_4_in_key_empty;
wire [127 : 0] expand_key2_128_4_out_key_data;
wire expand_key2_128_4_out_key_wr;
wire expand_key2_128_4_out_key_full;
	
// actor expand_key3_128_4
wire [127 : 0] fifo_small_expand_key3_128_4_in_key_data;
wire fifo_small_expand_key3_128_4_in_key_wr;
wire fifo_small_expand_key3_128_4_in_key_full;
wire [127 : 0] expand_key3_128_4_in_key_data;
wire expand_key3_128_4_in_key_rd;
wire expand_key3_128_4_in_key_empty;
wire [127 : 0] expand_key3_128_4_out_key_data;
wire expand_key3_128_4_out_key_wr;
wire expand_key3_128_4_out_key_full;
	
// actor expand_key0_128_5
wire [127 : 0] fifo_small_expand_key0_128_5_in_key_data;
wire fifo_small_expand_key0_128_5_in_key_wr;
wire fifo_small_expand_key0_128_5_in_key_full;
wire [127 : 0] expand_key0_128_5_in_key_data;
wire expand_key0_128_5_in_key_rd;
wire expand_key0_128_5_in_key_empty;
wire [7 : 0] fifo_small_expand_key0_128_5_in_rc_data;
wire fifo_small_expand_key0_128_5_in_rc_wr;
wire fifo_small_expand_key0_128_5_in_rc_full;
wire [7 : 0] expand_key0_128_5_in_rc_data;
wire expand_key0_128_5_in_rc_rd;
wire expand_key0_128_5_in_rc_empty;
wire [127 : 0] expand_key0_128_5_out_key_data;
wire expand_key0_128_5_out_key_wr;
wire expand_key0_128_5_out_key_full;
	
// actor expand_key1_128_5
wire [127 : 0] fifo_small_expand_key1_128_5_in_key_data;
wire fifo_small_expand_key1_128_5_in_key_wr;
wire fifo_small_expand_key1_128_5_in_key_full;
wire [127 : 0] expand_key1_128_5_in_key_data;
wire expand_key1_128_5_in_key_rd;
wire expand_key1_128_5_in_key_empty;
wire [127 : 0] expand_key1_128_5_out_key_data;
wire expand_key1_128_5_out_key_wr;
wire expand_key1_128_5_out_key_full;
	
// actor expand_key2_128_5
wire [127 : 0] fifo_small_expand_key2_128_5_in_key_data;
wire fifo_small_expand_key2_128_5_in_key_wr;
wire fifo_small_expand_key2_128_5_in_key_full;
wire [127 : 0] expand_key2_128_5_in_key_data;
wire expand_key2_128_5_in_key_rd;
wire expand_key2_128_5_in_key_empty;
wire [127 : 0] expand_key2_128_5_out_key_data;
wire expand_key2_128_5_out_key_wr;
wire expand_key2_128_5_out_key_full;
	
// actor expand_key3_128_5
wire [127 : 0] fifo_small_expand_key3_128_5_in_key_data;
wire fifo_small_expand_key3_128_5_in_key_wr;
wire fifo_small_expand_key3_128_5_in_key_full;
wire [127 : 0] expand_key3_128_5_in_key_data;
wire expand_key3_128_5_in_key_rd;
wire expand_key3_128_5_in_key_empty;
wire [127 : 0] expand_key3_128_5_out_key_data;
wire expand_key3_128_5_out_key_wr;
wire expand_key3_128_5_out_key_full;
	
// actor expand_key0_128_6
wire [127 : 0] fifo_small_expand_key0_128_6_in_key_data;
wire fifo_small_expand_key0_128_6_in_key_wr;
wire fifo_small_expand_key0_128_6_in_key_full;
wire [127 : 0] expand_key0_128_6_in_key_data;
wire expand_key0_128_6_in_key_rd;
wire expand_key0_128_6_in_key_empty;
wire [7 : 0] fifo_small_expand_key0_128_6_in_rc_data;
wire fifo_small_expand_key0_128_6_in_rc_wr;
wire fifo_small_expand_key0_128_6_in_rc_full;
wire [7 : 0] expand_key0_128_6_in_rc_data;
wire expand_key0_128_6_in_rc_rd;
wire expand_key0_128_6_in_rc_empty;
wire [127 : 0] expand_key0_128_6_out_key_data;
wire expand_key0_128_6_out_key_wr;
wire expand_key0_128_6_out_key_full;
	
// actor expand_key1_128_6
wire [127 : 0] fifo_small_expand_key1_128_6_in_key_data;
wire fifo_small_expand_key1_128_6_in_key_wr;
wire fifo_small_expand_key1_128_6_in_key_full;
wire [127 : 0] expand_key1_128_6_in_key_data;
wire expand_key1_128_6_in_key_rd;
wire expand_key1_128_6_in_key_empty;
wire [127 : 0] expand_key1_128_6_out_key_data;
wire expand_key1_128_6_out_key_wr;
wire expand_key1_128_6_out_key_full;
	
// actor expand_key2_128_6
wire [127 : 0] fifo_small_expand_key2_128_6_in_key_data;
wire fifo_small_expand_key2_128_6_in_key_wr;
wire fifo_small_expand_key2_128_6_in_key_full;
wire [127 : 0] expand_key2_128_6_in_key_data;
wire expand_key2_128_6_in_key_rd;
wire expand_key2_128_6_in_key_empty;
wire [127 : 0] expand_key2_128_6_out_key_data;
wire expand_key2_128_6_out_key_wr;
wire expand_key2_128_6_out_key_full;
	
// actor expand_key3_128_6
wire [127 : 0] fifo_small_expand_key3_128_6_in_key_data;
wire fifo_small_expand_key3_128_6_in_key_wr;
wire fifo_small_expand_key3_128_6_in_key_full;
wire [127 : 0] expand_key3_128_6_in_key_data;
wire expand_key3_128_6_in_key_rd;
wire expand_key3_128_6_in_key_empty;
wire [127 : 0] expand_key3_128_6_out_key_data;
wire expand_key3_128_6_out_key_wr;
wire expand_key3_128_6_out_key_full;
	
// actor expand_key0_128_7
wire [127 : 0] fifo_small_expand_key0_128_7_in_key_data;
wire fifo_small_expand_key0_128_7_in_key_wr;
wire fifo_small_expand_key0_128_7_in_key_full;
wire [127 : 0] expand_key0_128_7_in_key_data;
wire expand_key0_128_7_in_key_rd;
wire expand_key0_128_7_in_key_empty;
wire [7 : 0] fifo_small_expand_key0_128_7_in_rc_data;
wire fifo_small_expand_key0_128_7_in_rc_wr;
wire fifo_small_expand_key0_128_7_in_rc_full;
wire [7 : 0] expand_key0_128_7_in_rc_data;
wire expand_key0_128_7_in_rc_rd;
wire expand_key0_128_7_in_rc_empty;
wire [127 : 0] expand_key0_128_7_out_key_data;
wire expand_key0_128_7_out_key_wr;
wire expand_key0_128_7_out_key_full;
	
// actor expand_key1_128_7
wire [127 : 0] fifo_small_expand_key1_128_7_in_key_data;
wire fifo_small_expand_key1_128_7_in_key_wr;
wire fifo_small_expand_key1_128_7_in_key_full;
wire [127 : 0] expand_key1_128_7_in_key_data;
wire expand_key1_128_7_in_key_rd;
wire expand_key1_128_7_in_key_empty;
wire [127 : 0] expand_key1_128_7_out_key_data;
wire expand_key1_128_7_out_key_wr;
wire expand_key1_128_7_out_key_full;
	
// actor expand_key2_128_7
wire [127 : 0] fifo_small_expand_key2_128_7_in_key_data;
wire fifo_small_expand_key2_128_7_in_key_wr;
wire fifo_small_expand_key2_128_7_in_key_full;
wire [127 : 0] expand_key2_128_7_in_key_data;
wire expand_key2_128_7_in_key_rd;
wire expand_key2_128_7_in_key_empty;
wire [127 : 0] expand_key2_128_7_out_key_data;
wire expand_key2_128_7_out_key_wr;
wire expand_key2_128_7_out_key_full;
	
// actor expand_key3_128_7
wire [127 : 0] fifo_small_expand_key3_128_7_in_key_data;
wire fifo_small_expand_key3_128_7_in_key_wr;
wire fifo_small_expand_key3_128_7_in_key_full;
wire [127 : 0] expand_key3_128_7_in_key_data;
wire expand_key3_128_7_in_key_rd;
wire expand_key3_128_7_in_key_empty;
wire [127 : 0] expand_key3_128_7_out_key_data;
wire expand_key3_128_7_out_key_wr;
wire expand_key3_128_7_out_key_full;
	
// actor expand_key0_128_8
wire [127 : 0] fifo_small_expand_key0_128_8_in_key_data;
wire fifo_small_expand_key0_128_8_in_key_wr;
wire fifo_small_expand_key0_128_8_in_key_full;
wire [127 : 0] expand_key0_128_8_in_key_data;
wire expand_key0_128_8_in_key_rd;
wire expand_key0_128_8_in_key_empty;
wire [7 : 0] fifo_small_expand_key0_128_8_in_rc_data;
wire fifo_small_expand_key0_128_8_in_rc_wr;
wire fifo_small_expand_key0_128_8_in_rc_full;
wire [7 : 0] expand_key0_128_8_in_rc_data;
wire expand_key0_128_8_in_rc_rd;
wire expand_key0_128_8_in_rc_empty;
wire [127 : 0] expand_key0_128_8_out_key_data;
wire expand_key0_128_8_out_key_wr;
wire expand_key0_128_8_out_key_full;
	
// actor expand_key1_128_8
wire [127 : 0] fifo_small_expand_key1_128_8_in_key_data;
wire fifo_small_expand_key1_128_8_in_key_wr;
wire fifo_small_expand_key1_128_8_in_key_full;
wire [127 : 0] expand_key1_128_8_in_key_data;
wire expand_key1_128_8_in_key_rd;
wire expand_key1_128_8_in_key_empty;
wire [127 : 0] expand_key1_128_8_out_key_data;
wire expand_key1_128_8_out_key_wr;
wire expand_key1_128_8_out_key_full;
	
// actor expand_key2_128_8
wire [127 : 0] fifo_small_expand_key2_128_8_in_key_data;
wire fifo_small_expand_key2_128_8_in_key_wr;
wire fifo_small_expand_key2_128_8_in_key_full;
wire [127 : 0] expand_key2_128_8_in_key_data;
wire expand_key2_128_8_in_key_rd;
wire expand_key2_128_8_in_key_empty;
wire [127 : 0] expand_key2_128_8_out_key_data;
wire expand_key2_128_8_out_key_wr;
wire expand_key2_128_8_out_key_full;
	
// actor expand_key3_128_8
wire [127 : 0] fifo_small_expand_key3_128_8_in_key_data;
wire fifo_small_expand_key3_128_8_in_key_wr;
wire fifo_small_expand_key3_128_8_in_key_full;
wire [127 : 0] expand_key3_128_8_in_key_data;
wire expand_key3_128_8_in_key_rd;
wire expand_key3_128_8_in_key_empty;
wire [127 : 0] expand_key3_128_8_out_key_data;
wire expand_key3_128_8_out_key_wr;
wire expand_key3_128_8_out_key_full;
	
// actor sub_bytes_9
wire [127 : 0] fifo_small_sub_bytes_9_in_state_data;
wire fifo_small_sub_bytes_9_in_state_wr;
wire fifo_small_sub_bytes_9_in_state_full;
wire [127 : 0] sub_bytes_9_in_state_data;
wire sub_bytes_9_in_state_rd;
wire sub_bytes_9_in_state_empty;
wire [127 : 0] sub_bytes_9_out_state_data;
wire sub_bytes_9_out_state_wr;
wire sub_bytes_9_out_state_full;
	
// actor shift_rows_9
wire [127 : 0] fifo_small_shift_rows_9_in_state_data;
wire fifo_small_shift_rows_9_in_state_wr;
wire fifo_small_shift_rows_9_in_state_full;
wire [127 : 0] shift_rows_9_in_state_data;
wire shift_rows_9_in_state_rd;
wire shift_rows_9_in_state_empty;
wire [127 : 0] shift_rows_9_out_state_data;
wire shift_rows_9_out_state_wr;
wire shift_rows_9_out_state_full;
	
// actor mix_cols_8
wire [127 : 0] fifo_small_mix_cols_8_in_state_data;
wire fifo_small_mix_cols_8_in_state_wr;
wire fifo_small_mix_cols_8_in_state_full;
wire [127 : 0] mix_cols_8_in_state_data;
wire mix_cols_8_in_state_rd;
wire mix_cols_8_in_state_empty;
wire [127 : 0] mix_cols_8_out_state_data;
wire mix_cols_8_out_state_wr;
wire mix_cols_8_out_state_full;
	
// actor add_round_key_10
wire [127 : 0] fifo_small_add_round_key_10_in_state_data;
wire fifo_small_add_round_key_10_in_state_wr;
wire fifo_small_add_round_key_10_in_state_full;
wire [127 : 0] add_round_key_10_in_state_data;
wire add_round_key_10_in_state_rd;
wire add_round_key_10_in_state_empty;
wire [127 : 0] fifo_small_add_round_key_10_round_key_data;
wire fifo_small_add_round_key_10_round_key_wr;
wire fifo_small_add_round_key_10_round_key_full;
wire [127 : 0] add_round_key_10_round_key_data;
wire add_round_key_10_round_key_rd;
wire add_round_key_10_round_key_empty;
wire [127 : 0] add_round_key_10_out_state_data;
wire add_round_key_10_out_state_wr;
wire add_round_key_10_out_state_full;
	
// actor expand_key0_128_9
wire [127 : 0] fifo_small_expand_key0_128_9_in_key_data;
wire fifo_small_expand_key0_128_9_in_key_wr;
wire fifo_small_expand_key0_128_9_in_key_full;
wire [127 : 0] expand_key0_128_9_in_key_data;
wire expand_key0_128_9_in_key_rd;
wire expand_key0_128_9_in_key_empty;
wire [7 : 0] fifo_small_expand_key0_128_9_in_rc_data;
wire fifo_small_expand_key0_128_9_in_rc_wr;
wire fifo_small_expand_key0_128_9_in_rc_full;
wire [7 : 0] expand_key0_128_9_in_rc_data;
wire expand_key0_128_9_in_rc_rd;
wire expand_key0_128_9_in_rc_empty;
wire [127 : 0] expand_key0_128_9_out_key_data;
wire expand_key0_128_9_out_key_wr;
wire expand_key0_128_9_out_key_full;
	
// actor expand_key1_128_9
wire [127 : 0] fifo_small_expand_key1_128_9_in_key_data;
wire fifo_small_expand_key1_128_9_in_key_wr;
wire fifo_small_expand_key1_128_9_in_key_full;
wire [127 : 0] expand_key1_128_9_in_key_data;
wire expand_key1_128_9_in_key_rd;
wire expand_key1_128_9_in_key_empty;
wire [127 : 0] expand_key1_128_9_out_key_data;
wire expand_key1_128_9_out_key_wr;
wire expand_key1_128_9_out_key_full;
	
// actor expand_key2_128_9
wire [127 : 0] fifo_small_expand_key2_128_9_in_key_data;
wire fifo_small_expand_key2_128_9_in_key_wr;
wire fifo_small_expand_key2_128_9_in_key_full;
wire [127 : 0] expand_key2_128_9_in_key_data;
wire expand_key2_128_9_in_key_rd;
wire expand_key2_128_9_in_key_empty;
wire [127 : 0] expand_key2_128_9_out_key_data;
wire expand_key2_128_9_out_key_wr;
wire expand_key2_128_9_out_key_full;
	
// actor expand_key3_128_9
wire [127 : 0] fifo_small_expand_key3_128_9_in_key_data;
wire fifo_small_expand_key3_128_9_in_key_wr;
wire fifo_small_expand_key3_128_9_in_key_full;
wire [127 : 0] expand_key3_128_9_in_key_data;
wire expand_key3_128_9_in_key_rd;
wire expand_key3_128_9_in_key_empty;
wire [127 : 0] expand_key3_128_9_out_key_data;
wire expand_key3_128_9_out_key_wr;
wire expand_key3_128_9_out_key_full;
// ----------------------------------------------------------------------------

// body
// ----------------------------------------------------------------------------



// fifo_small_add_round_key_0_in_state
fifo_small #(
	.depth(64),
	.size(128)
) fifo_small_add_round_key_0_in_state(
	.datain(fifo_small_add_round_key_0_in_state_data),
	.dataout(add_round_key_0_in_state_data),
	.enr(add_round_key_0_in_state_rd),
	.enw(fifo_small_add_round_key_0_in_state_wr),
	.empty(add_round_key_0_in_state_empty),
	.full(fifo_small_add_round_key_0_in_state_full),
	
	// System Signal(s)
	.clk(clock),
	.rst(reset)
);
// fifo_small_add_round_key_0_round_key
fifo_small #(
	.depth(64),
	.size(128)
) fifo_small_add_round_key_0_round_key(
	.datain(fifo_small_add_round_key_0_round_key_data),
	.dataout(add_round_key_0_round_key_data),
	.enr(add_round_key_0_round_key_rd),
	.enw(fifo_small_add_round_key_0_round_key_wr),
	.empty(add_round_key_0_round_key_empty),
	.full(fifo_small_add_round_key_0_round_key_full),
	
	// System Signal(s)
	.clk(clock),
	.rst(reset)
);

// actor add_round_key_0
add_round_key actor_add_round_key_0 (
	// Input Signal(s)
	.in_state(add_round_key_0_in_state_data),
	.in_state_rd(add_round_key_0_in_state_rd),
	.in_state_empty(add_round_key_0_in_state_empty),
	.round_key(add_round_key_0_round_key_data),
	.round_key_rd(add_round_key_0_round_key_rd),
	.round_key_empty(add_round_key_0_round_key_empty)
	,
	
	// Output Signal(s)
	.out_state(add_round_key_0_out_state_data),
	.out_state_wr(add_round_key_0_out_state_wr),
	.out_state_full(add_round_key_0_out_state_full)
		,
	
	// System Signal(s)
	.clock(clock),
	.reset(reset)
);


// fifo_small_sub_bytes_0_in_state
fifo_small #(
	.depth(64),
	.size(128)
) fifo_small_sub_bytes_0_in_state(
	.datain(fifo_small_sub_bytes_0_in_state_data),
	.dataout(sub_bytes_0_in_state_data),
	.enr(sub_bytes_0_in_state_rd),
	.enw(fifo_small_sub_bytes_0_in_state_wr),
	.empty(sub_bytes_0_in_state_empty),
	.full(fifo_small_sub_bytes_0_in_state_full),
	
	// System Signal(s)
	.clk(clock),
	.rst(reset)
);

// actor sub_bytes_0
sub_bytes actor_sub_bytes_0 (
	// Input Signal(s)
	.in_state(sub_bytes_0_in_state_data),
	.in_state_rd(sub_bytes_0_in_state_rd),
	.in_state_empty(sub_bytes_0_in_state_empty)
	,
	
	// Output Signal(s)
	.out_state(sub_bytes_0_out_state_data),
	.out_state_wr(sub_bytes_0_out_state_wr),
	.out_state_full(sub_bytes_0_out_state_full)
		,
	
	// System Signal(s)
	.clock(clock),
	.reset(reset)
);


// fifo_small_shift_rows_0_in_state
fifo_small #(
	.depth(64),
	.size(128)
) fifo_small_shift_rows_0_in_state(
	.datain(fifo_small_shift_rows_0_in_state_data),
	.dataout(shift_rows_0_in_state_data),
	.enr(shift_rows_0_in_state_rd),
	.enw(fifo_small_shift_rows_0_in_state_wr),
	.empty(shift_rows_0_in_state_empty),
	.full(fifo_small_shift_rows_0_in_state_full),
	
	// System Signal(s)
	.clk(clock),
	.rst(reset)
);

// actor shift_rows_0
shift_rows actor_shift_rows_0 (
	// Input Signal(s)
	.in_state(shift_rows_0_in_state_data),
	.in_state_rd(shift_rows_0_in_state_rd),
	.in_state_empty(shift_rows_0_in_state_empty)
	,
	
	// Output Signal(s)
	.out_state(shift_rows_0_out_state_data),
	.out_state_wr(shift_rows_0_out_state_wr),
	.out_state_full(shift_rows_0_out_state_full)
		,
	
	// System Signal(s)
	.clock(clock),
	.reset(reset)
);


// fifo_small_add_round_key_1_in_state
fifo_small #(
	.depth(64),
	.size(128)
) fifo_small_add_round_key_1_in_state(
	.datain(fifo_small_add_round_key_1_in_state_data),
	.dataout(add_round_key_1_in_state_data),
	.enr(add_round_key_1_in_state_rd),
	.enw(fifo_small_add_round_key_1_in_state_wr),
	.empty(add_round_key_1_in_state_empty),
	.full(fifo_small_add_round_key_1_in_state_full),
	
	// System Signal(s)
	.clk(clock),
	.rst(reset)
);
// fifo_small_add_round_key_1_round_key
fifo_small #(
	.depth(64),
	.size(128)
) fifo_small_add_round_key_1_round_key(
	.datain(fifo_small_add_round_key_1_round_key_data),
	.dataout(add_round_key_1_round_key_data),
	.enr(add_round_key_1_round_key_rd),
	.enw(fifo_small_add_round_key_1_round_key_wr),
	.empty(add_round_key_1_round_key_empty),
	.full(fifo_small_add_round_key_1_round_key_full),
	
	// System Signal(s)
	.clk(clock),
	.rst(reset)
);

// actor add_round_key_1
add_round_key actor_add_round_key_1 (
	// Input Signal(s)
	.in_state(add_round_key_1_in_state_data),
	.in_state_rd(add_round_key_1_in_state_rd),
	.in_state_empty(add_round_key_1_in_state_empty),
	.round_key(add_round_key_1_round_key_data),
	.round_key_rd(add_round_key_1_round_key_rd),
	.round_key_empty(add_round_key_1_round_key_empty)
	,
	
	// Output Signal(s)
	.out_state(add_round_key_1_out_state_data),
	.out_state_wr(add_round_key_1_out_state_wr),
	.out_state_full(add_round_key_1_out_state_full)
		,
	
	// System Signal(s)
	.clock(clock),
	.reset(reset)
);


// fifo_small_read8x16_0_in_token
fifo_small #(
	.depth(64),
	.size(8)
) fifo_small_read8x16_0_in_token(
	.datain(fifo_small_read8x16_0_in_token_data),
	.dataout(read8x16_0_in_token_data),
	.enr(read8x16_0_in_token_rd),
	.enw(fifo_small_read8x16_0_in_token_wr),
	.empty(read8x16_0_in_token_empty),
	.full(fifo_small_read8x16_0_in_token_full),
	
	// System Signal(s)
	.clk(clock),
	.rst(reset)
);

// actor read8x16_0
read8x16 actor_read8x16_0 (
	// Input Signal(s)
	.in_token(read8x16_0_in_token_data),
	.in_token_rd(read8x16_0_in_token_rd),
	.in_token_empty(read8x16_0_in_token_empty)
	,
	
	// Output Signal(s)
	.out_token(read8x16_0_out_token_data),
	.out_token_wr(read8x16_0_out_token_wr),
	.out_token_full(read8x16_0_out_token_full)
		,
	
	// System Signal(s)
	.clock(clock),
	.reset(reset)
);


// fifo_small_read8x16_1_in_token
fifo_small #(
	.depth(64),
	.size(8)
) fifo_small_read8x16_1_in_token(
	.datain(fifo_small_read8x16_1_in_token_data),
	.dataout(read8x16_1_in_token_data),
	.enr(read8x16_1_in_token_rd),
	.enw(fifo_small_read8x16_1_in_token_wr),
	.empty(read8x16_1_in_token_empty),
	.full(fifo_small_read8x16_1_in_token_full),
	
	// System Signal(s)
	.clk(clock),
	.rst(reset)
);

// actor read8x16_1
read8x16 actor_read8x16_1 (
	// Input Signal(s)
	.in_token(read8x16_1_in_token_data),
	.in_token_rd(read8x16_1_in_token_rd),
	.in_token_empty(read8x16_1_in_token_empty)
	,
	
	// Output Signal(s)
	.out_token(read8x16_1_out_token_data),
	.out_token_wr(read8x16_1_out_token_wr),
	.out_token_full(read8x16_1_out_token_full)
		,
	
	// System Signal(s)
	.clock(clock),
	.reset(reset)
);


// fifo_small_write16x8_0_in_token
fifo_small #(
	.depth(64),
	.size(128)
) fifo_small_write16x8_0_in_token(
	.datain(fifo_small_write16x8_0_in_token_data),
	.dataout(write16x8_0_in_token_data),
	.enr(write16x8_0_in_token_rd),
	.enw(fifo_small_write16x8_0_in_token_wr),
	.empty(write16x8_0_in_token_empty),
	.full(fifo_small_write16x8_0_in_token_full),
	
	// System Signal(s)
	.clk(clock),
	.rst(reset)
);

// actor write16x8_0
write16x8 actor_write16x8_0 (
	// Input Signal(s)
	.in_token(write16x8_0_in_token_data),
	.in_token_rd(write16x8_0_in_token_rd),
	.in_token_empty(write16x8_0_in_token_empty)
	,
	
	// Output Signal(s)
	.out_token(write16x8_0_out_token_data),
	.out_token_wr(write16x8_0_out_token_wr),
	.out_token_full(write16x8_0_out_token_full)
		,
	
	// System Signal(s)
	.clock(clock),
	.reset(reset)
);


// fifo_small_sub_bytes_1_in_state
fifo_small #(
	.depth(64),
	.size(128)
) fifo_small_sub_bytes_1_in_state(
	.datain(fifo_small_sub_bytes_1_in_state_data),
	.dataout(sub_bytes_1_in_state_data),
	.enr(sub_bytes_1_in_state_rd),
	.enw(fifo_small_sub_bytes_1_in_state_wr),
	.empty(sub_bytes_1_in_state_empty),
	.full(fifo_small_sub_bytes_1_in_state_full),
	
	// System Signal(s)
	.clk(clock),
	.rst(reset)
);

// actor sub_bytes_1
sub_bytes actor_sub_bytes_1 (
	// Input Signal(s)
	.in_state(sub_bytes_1_in_state_data),
	.in_state_rd(sub_bytes_1_in_state_rd),
	.in_state_empty(sub_bytes_1_in_state_empty)
	,
	
	// Output Signal(s)
	.out_state(sub_bytes_1_out_state_data),
	.out_state_wr(sub_bytes_1_out_state_wr),
	.out_state_full(sub_bytes_1_out_state_full)
		,
	
	// System Signal(s)
	.clock(clock),
	.reset(reset)
);


// fifo_small_shift_rows_1_in_state
fifo_small #(
	.depth(64),
	.size(128)
) fifo_small_shift_rows_1_in_state(
	.datain(fifo_small_shift_rows_1_in_state_data),
	.dataout(shift_rows_1_in_state_data),
	.enr(shift_rows_1_in_state_rd),
	.enw(fifo_small_shift_rows_1_in_state_wr),
	.empty(shift_rows_1_in_state_empty),
	.full(fifo_small_shift_rows_1_in_state_full),
	
	// System Signal(s)
	.clk(clock),
	.rst(reset)
);

// actor shift_rows_1
shift_rows actor_shift_rows_1 (
	// Input Signal(s)
	.in_state(shift_rows_1_in_state_data),
	.in_state_rd(shift_rows_1_in_state_rd),
	.in_state_empty(shift_rows_1_in_state_empty)
	,
	
	// Output Signal(s)
	.out_state(shift_rows_1_out_state_data),
	.out_state_wr(shift_rows_1_out_state_wr),
	.out_state_full(shift_rows_1_out_state_full)
		,
	
	// System Signal(s)
	.clock(clock),
	.reset(reset)
);


// fifo_small_mix_cols_0_in_state
fifo_small #(
	.depth(64),
	.size(128)
) fifo_small_mix_cols_0_in_state(
	.datain(fifo_small_mix_cols_0_in_state_data),
	.dataout(mix_cols_0_in_state_data),
	.enr(mix_cols_0_in_state_rd),
	.enw(fifo_small_mix_cols_0_in_state_wr),
	.empty(mix_cols_0_in_state_empty),
	.full(fifo_small_mix_cols_0_in_state_full),
	
	// System Signal(s)
	.clk(clock),
	.rst(reset)
);

// actor mix_cols_0
mix_cols actor_mix_cols_0 (
	// Input Signal(s)
	.in_state(mix_cols_0_in_state_data),
	.in_state_rd(mix_cols_0_in_state_rd),
	.in_state_empty(mix_cols_0_in_state_empty)
	,
	
	// Output Signal(s)
	.out_state(mix_cols_0_out_state_data),
	.out_state_wr(mix_cols_0_out_state_wr),
	.out_state_full(mix_cols_0_out_state_full)
		,
	
	// System Signal(s)
	.clock(clock),
	.reset(reset)
);


// fifo_small_add_round_key_2_in_state
fifo_small #(
	.depth(64),
	.size(128)
) fifo_small_add_round_key_2_in_state(
	.datain(fifo_small_add_round_key_2_in_state_data),
	.dataout(add_round_key_2_in_state_data),
	.enr(add_round_key_2_in_state_rd),
	.enw(fifo_small_add_round_key_2_in_state_wr),
	.empty(add_round_key_2_in_state_empty),
	.full(fifo_small_add_round_key_2_in_state_full),
	
	// System Signal(s)
	.clk(clock),
	.rst(reset)
);
// fifo_small_add_round_key_2_round_key
fifo_small #(
	.depth(64),
	.size(128)
) fifo_small_add_round_key_2_round_key(
	.datain(fifo_small_add_round_key_2_round_key_data),
	.dataout(add_round_key_2_round_key_data),
	.enr(add_round_key_2_round_key_rd),
	.enw(fifo_small_add_round_key_2_round_key_wr),
	.empty(add_round_key_2_round_key_empty),
	.full(fifo_small_add_round_key_2_round_key_full),
	
	// System Signal(s)
	.clk(clock),
	.rst(reset)
);

// actor add_round_key_2
add_round_key actor_add_round_key_2 (
	// Input Signal(s)
	.in_state(add_round_key_2_in_state_data),
	.in_state_rd(add_round_key_2_in_state_rd),
	.in_state_empty(add_round_key_2_in_state_empty),
	.round_key(add_round_key_2_round_key_data),
	.round_key_rd(add_round_key_2_round_key_rd),
	.round_key_empty(add_round_key_2_round_key_empty)
	,
	
	// Output Signal(s)
	.out_state(add_round_key_2_out_state_data),
	.out_state_wr(add_round_key_2_out_state_wr),
	.out_state_full(add_round_key_2_out_state_full)
		,
	
	// System Signal(s)
	.clock(clock),
	.reset(reset)
);


// fifo_small_sub_bytes_2_in_state
fifo_small #(
	.depth(64),
	.size(128)
) fifo_small_sub_bytes_2_in_state(
	.datain(fifo_small_sub_bytes_2_in_state_data),
	.dataout(sub_bytes_2_in_state_data),
	.enr(sub_bytes_2_in_state_rd),
	.enw(fifo_small_sub_bytes_2_in_state_wr),
	.empty(sub_bytes_2_in_state_empty),
	.full(fifo_small_sub_bytes_2_in_state_full),
	
	// System Signal(s)
	.clk(clock),
	.rst(reset)
);

// actor sub_bytes_2
sub_bytes actor_sub_bytes_2 (
	// Input Signal(s)
	.in_state(sub_bytes_2_in_state_data),
	.in_state_rd(sub_bytes_2_in_state_rd),
	.in_state_empty(sub_bytes_2_in_state_empty)
	,
	
	// Output Signal(s)
	.out_state(sub_bytes_2_out_state_data),
	.out_state_wr(sub_bytes_2_out_state_wr),
	.out_state_full(sub_bytes_2_out_state_full)
		,
	
	// System Signal(s)
	.clock(clock),
	.reset(reset)
);


// fifo_small_shift_rows_2_in_state
fifo_small #(
	.depth(64),
	.size(128)
) fifo_small_shift_rows_2_in_state(
	.datain(fifo_small_shift_rows_2_in_state_data),
	.dataout(shift_rows_2_in_state_data),
	.enr(shift_rows_2_in_state_rd),
	.enw(fifo_small_shift_rows_2_in_state_wr),
	.empty(shift_rows_2_in_state_empty),
	.full(fifo_small_shift_rows_2_in_state_full),
	
	// System Signal(s)
	.clk(clock),
	.rst(reset)
);

// actor shift_rows_2
shift_rows actor_shift_rows_2 (
	// Input Signal(s)
	.in_state(shift_rows_2_in_state_data),
	.in_state_rd(shift_rows_2_in_state_rd),
	.in_state_empty(shift_rows_2_in_state_empty)
	,
	
	// Output Signal(s)
	.out_state(shift_rows_2_out_state_data),
	.out_state_wr(shift_rows_2_out_state_wr),
	.out_state_full(shift_rows_2_out_state_full)
		,
	
	// System Signal(s)
	.clock(clock),
	.reset(reset)
);


// fifo_small_mix_cols_1_in_state
fifo_small #(
	.depth(64),
	.size(128)
) fifo_small_mix_cols_1_in_state(
	.datain(fifo_small_mix_cols_1_in_state_data),
	.dataout(mix_cols_1_in_state_data),
	.enr(mix_cols_1_in_state_rd),
	.enw(fifo_small_mix_cols_1_in_state_wr),
	.empty(mix_cols_1_in_state_empty),
	.full(fifo_small_mix_cols_1_in_state_full),
	
	// System Signal(s)
	.clk(clock),
	.rst(reset)
);

// actor mix_cols_1
mix_cols actor_mix_cols_1 (
	// Input Signal(s)
	.in_state(mix_cols_1_in_state_data),
	.in_state_rd(mix_cols_1_in_state_rd),
	.in_state_empty(mix_cols_1_in_state_empty)
	,
	
	// Output Signal(s)
	.out_state(mix_cols_1_out_state_data),
	.out_state_wr(mix_cols_1_out_state_wr),
	.out_state_full(mix_cols_1_out_state_full)
		,
	
	// System Signal(s)
	.clock(clock),
	.reset(reset)
);


// fifo_small_add_round_key_3_in_state
fifo_small #(
	.depth(64),
	.size(128)
) fifo_small_add_round_key_3_in_state(
	.datain(fifo_small_add_round_key_3_in_state_data),
	.dataout(add_round_key_3_in_state_data),
	.enr(add_round_key_3_in_state_rd),
	.enw(fifo_small_add_round_key_3_in_state_wr),
	.empty(add_round_key_3_in_state_empty),
	.full(fifo_small_add_round_key_3_in_state_full),
	
	// System Signal(s)
	.clk(clock),
	.rst(reset)
);
// fifo_small_add_round_key_3_round_key
fifo_small #(
	.depth(64),
	.size(128)
) fifo_small_add_round_key_3_round_key(
	.datain(fifo_small_add_round_key_3_round_key_data),
	.dataout(add_round_key_3_round_key_data),
	.enr(add_round_key_3_round_key_rd),
	.enw(fifo_small_add_round_key_3_round_key_wr),
	.empty(add_round_key_3_round_key_empty),
	.full(fifo_small_add_round_key_3_round_key_full),
	
	// System Signal(s)
	.clk(clock),
	.rst(reset)
);

// actor add_round_key_3
add_round_key actor_add_round_key_3 (
	// Input Signal(s)
	.in_state(add_round_key_3_in_state_data),
	.in_state_rd(add_round_key_3_in_state_rd),
	.in_state_empty(add_round_key_3_in_state_empty),
	.round_key(add_round_key_3_round_key_data),
	.round_key_rd(add_round_key_3_round_key_rd),
	.round_key_empty(add_round_key_3_round_key_empty)
	,
	
	// Output Signal(s)
	.out_state(add_round_key_3_out_state_data),
	.out_state_wr(add_round_key_3_out_state_wr),
	.out_state_full(add_round_key_3_out_state_full)
		,
	
	// System Signal(s)
	.clock(clock),
	.reset(reset)
);


// fifo_small_sub_bytes_3_in_state
fifo_small #(
	.depth(64),
	.size(128)
) fifo_small_sub_bytes_3_in_state(
	.datain(fifo_small_sub_bytes_3_in_state_data),
	.dataout(sub_bytes_3_in_state_data),
	.enr(sub_bytes_3_in_state_rd),
	.enw(fifo_small_sub_bytes_3_in_state_wr),
	.empty(sub_bytes_3_in_state_empty),
	.full(fifo_small_sub_bytes_3_in_state_full),
	
	// System Signal(s)
	.clk(clock),
	.rst(reset)
);

// actor sub_bytes_3
sub_bytes actor_sub_bytes_3 (
	// Input Signal(s)
	.in_state(sub_bytes_3_in_state_data),
	.in_state_rd(sub_bytes_3_in_state_rd),
	.in_state_empty(sub_bytes_3_in_state_empty)
	,
	
	// Output Signal(s)
	.out_state(sub_bytes_3_out_state_data),
	.out_state_wr(sub_bytes_3_out_state_wr),
	.out_state_full(sub_bytes_3_out_state_full)
		,
	
	// System Signal(s)
	.clock(clock),
	.reset(reset)
);


// fifo_small_shift_rows_3_in_state
fifo_small #(
	.depth(64),
	.size(128)
) fifo_small_shift_rows_3_in_state(
	.datain(fifo_small_shift_rows_3_in_state_data),
	.dataout(shift_rows_3_in_state_data),
	.enr(shift_rows_3_in_state_rd),
	.enw(fifo_small_shift_rows_3_in_state_wr),
	.empty(shift_rows_3_in_state_empty),
	.full(fifo_small_shift_rows_3_in_state_full),
	
	// System Signal(s)
	.clk(clock),
	.rst(reset)
);

// actor shift_rows_3
shift_rows actor_shift_rows_3 (
	// Input Signal(s)
	.in_state(shift_rows_3_in_state_data),
	.in_state_rd(shift_rows_3_in_state_rd),
	.in_state_empty(shift_rows_3_in_state_empty)
	,
	
	// Output Signal(s)
	.out_state(shift_rows_3_out_state_data),
	.out_state_wr(shift_rows_3_out_state_wr),
	.out_state_full(shift_rows_3_out_state_full)
		,
	
	// System Signal(s)
	.clock(clock),
	.reset(reset)
);


// fifo_small_mix_cols_2_in_state
fifo_small #(
	.depth(64),
	.size(128)
) fifo_small_mix_cols_2_in_state(
	.datain(fifo_small_mix_cols_2_in_state_data),
	.dataout(mix_cols_2_in_state_data),
	.enr(mix_cols_2_in_state_rd),
	.enw(fifo_small_mix_cols_2_in_state_wr),
	.empty(mix_cols_2_in_state_empty),
	.full(fifo_small_mix_cols_2_in_state_full),
	
	// System Signal(s)
	.clk(clock),
	.rst(reset)
);

// actor mix_cols_2
mix_cols actor_mix_cols_2 (
	// Input Signal(s)
	.in_state(mix_cols_2_in_state_data),
	.in_state_rd(mix_cols_2_in_state_rd),
	.in_state_empty(mix_cols_2_in_state_empty)
	,
	
	// Output Signal(s)
	.out_state(mix_cols_2_out_state_data),
	.out_state_wr(mix_cols_2_out_state_wr),
	.out_state_full(mix_cols_2_out_state_full)
		,
	
	// System Signal(s)
	.clock(clock),
	.reset(reset)
);


// fifo_small_add_round_key_4_in_state
fifo_small #(
	.depth(64),
	.size(128)
) fifo_small_add_round_key_4_in_state(
	.datain(fifo_small_add_round_key_4_in_state_data),
	.dataout(add_round_key_4_in_state_data),
	.enr(add_round_key_4_in_state_rd),
	.enw(fifo_small_add_round_key_4_in_state_wr),
	.empty(add_round_key_4_in_state_empty),
	.full(fifo_small_add_round_key_4_in_state_full),
	
	// System Signal(s)
	.clk(clock),
	.rst(reset)
);
// fifo_small_add_round_key_4_round_key
fifo_small #(
	.depth(64),
	.size(128)
) fifo_small_add_round_key_4_round_key(
	.datain(fifo_small_add_round_key_4_round_key_data),
	.dataout(add_round_key_4_round_key_data),
	.enr(add_round_key_4_round_key_rd),
	.enw(fifo_small_add_round_key_4_round_key_wr),
	.empty(add_round_key_4_round_key_empty),
	.full(fifo_small_add_round_key_4_round_key_full),
	
	// System Signal(s)
	.clk(clock),
	.rst(reset)
);

// actor add_round_key_4
add_round_key actor_add_round_key_4 (
	// Input Signal(s)
	.in_state(add_round_key_4_in_state_data),
	.in_state_rd(add_round_key_4_in_state_rd),
	.in_state_empty(add_round_key_4_in_state_empty),
	.round_key(add_round_key_4_round_key_data),
	.round_key_rd(add_round_key_4_round_key_rd),
	.round_key_empty(add_round_key_4_round_key_empty)
	,
	
	// Output Signal(s)
	.out_state(add_round_key_4_out_state_data),
	.out_state_wr(add_round_key_4_out_state_wr),
	.out_state_full(add_round_key_4_out_state_full)
		,
	
	// System Signal(s)
	.clock(clock),
	.reset(reset)
);


// fifo_small_sub_bytes_4_in_state
fifo_small #(
	.depth(64),
	.size(128)
) fifo_small_sub_bytes_4_in_state(
	.datain(fifo_small_sub_bytes_4_in_state_data),
	.dataout(sub_bytes_4_in_state_data),
	.enr(sub_bytes_4_in_state_rd),
	.enw(fifo_small_sub_bytes_4_in_state_wr),
	.empty(sub_bytes_4_in_state_empty),
	.full(fifo_small_sub_bytes_4_in_state_full),
	
	// System Signal(s)
	.clk(clock),
	.rst(reset)
);

// actor sub_bytes_4
sub_bytes actor_sub_bytes_4 (
	// Input Signal(s)
	.in_state(sub_bytes_4_in_state_data),
	.in_state_rd(sub_bytes_4_in_state_rd),
	.in_state_empty(sub_bytes_4_in_state_empty)
	,
	
	// Output Signal(s)
	.out_state(sub_bytes_4_out_state_data),
	.out_state_wr(sub_bytes_4_out_state_wr),
	.out_state_full(sub_bytes_4_out_state_full)
		,
	
	// System Signal(s)
	.clock(clock),
	.reset(reset)
);


// fifo_small_shift_rows_4_in_state
fifo_small #(
	.depth(64),
	.size(128)
) fifo_small_shift_rows_4_in_state(
	.datain(fifo_small_shift_rows_4_in_state_data),
	.dataout(shift_rows_4_in_state_data),
	.enr(shift_rows_4_in_state_rd),
	.enw(fifo_small_shift_rows_4_in_state_wr),
	.empty(shift_rows_4_in_state_empty),
	.full(fifo_small_shift_rows_4_in_state_full),
	
	// System Signal(s)
	.clk(clock),
	.rst(reset)
);

// actor shift_rows_4
shift_rows actor_shift_rows_4 (
	// Input Signal(s)
	.in_state(shift_rows_4_in_state_data),
	.in_state_rd(shift_rows_4_in_state_rd),
	.in_state_empty(shift_rows_4_in_state_empty)
	,
	
	// Output Signal(s)
	.out_state(shift_rows_4_out_state_data),
	.out_state_wr(shift_rows_4_out_state_wr),
	.out_state_full(shift_rows_4_out_state_full)
		,
	
	// System Signal(s)
	.clock(clock),
	.reset(reset)
);


// fifo_small_mix_cols_3_in_state
fifo_small #(
	.depth(64),
	.size(128)
) fifo_small_mix_cols_3_in_state(
	.datain(fifo_small_mix_cols_3_in_state_data),
	.dataout(mix_cols_3_in_state_data),
	.enr(mix_cols_3_in_state_rd),
	.enw(fifo_small_mix_cols_3_in_state_wr),
	.empty(mix_cols_3_in_state_empty),
	.full(fifo_small_mix_cols_3_in_state_full),
	
	// System Signal(s)
	.clk(clock),
	.rst(reset)
);

// actor mix_cols_3
mix_cols actor_mix_cols_3 (
	// Input Signal(s)
	.in_state(mix_cols_3_in_state_data),
	.in_state_rd(mix_cols_3_in_state_rd),
	.in_state_empty(mix_cols_3_in_state_empty)
	,
	
	// Output Signal(s)
	.out_state(mix_cols_3_out_state_data),
	.out_state_wr(mix_cols_3_out_state_wr),
	.out_state_full(mix_cols_3_out_state_full)
		,
	
	// System Signal(s)
	.clock(clock),
	.reset(reset)
);


// fifo_small_add_round_key_5_in_state
fifo_small #(
	.depth(64),
	.size(128)
) fifo_small_add_round_key_5_in_state(
	.datain(fifo_small_add_round_key_5_in_state_data),
	.dataout(add_round_key_5_in_state_data),
	.enr(add_round_key_5_in_state_rd),
	.enw(fifo_small_add_round_key_5_in_state_wr),
	.empty(add_round_key_5_in_state_empty),
	.full(fifo_small_add_round_key_5_in_state_full),
	
	// System Signal(s)
	.clk(clock),
	.rst(reset)
);
// fifo_small_add_round_key_5_round_key
fifo_small #(
	.depth(64),
	.size(128)
) fifo_small_add_round_key_5_round_key(
	.datain(fifo_small_add_round_key_5_round_key_data),
	.dataout(add_round_key_5_round_key_data),
	.enr(add_round_key_5_round_key_rd),
	.enw(fifo_small_add_round_key_5_round_key_wr),
	.empty(add_round_key_5_round_key_empty),
	.full(fifo_small_add_round_key_5_round_key_full),
	
	// System Signal(s)
	.clk(clock),
	.rst(reset)
);

// actor add_round_key_5
add_round_key actor_add_round_key_5 (
	// Input Signal(s)
	.in_state(add_round_key_5_in_state_data),
	.in_state_rd(add_round_key_5_in_state_rd),
	.in_state_empty(add_round_key_5_in_state_empty),
	.round_key(add_round_key_5_round_key_data),
	.round_key_rd(add_round_key_5_round_key_rd),
	.round_key_empty(add_round_key_5_round_key_empty)
	,
	
	// Output Signal(s)
	.out_state(add_round_key_5_out_state_data),
	.out_state_wr(add_round_key_5_out_state_wr),
	.out_state_full(add_round_key_5_out_state_full)
		,
	
	// System Signal(s)
	.clock(clock),
	.reset(reset)
);


// fifo_small_sub_bytes_5_in_state
fifo_small #(
	.depth(64),
	.size(128)
) fifo_small_sub_bytes_5_in_state(
	.datain(fifo_small_sub_bytes_5_in_state_data),
	.dataout(sub_bytes_5_in_state_data),
	.enr(sub_bytes_5_in_state_rd),
	.enw(fifo_small_sub_bytes_5_in_state_wr),
	.empty(sub_bytes_5_in_state_empty),
	.full(fifo_small_sub_bytes_5_in_state_full),
	
	// System Signal(s)
	.clk(clock),
	.rst(reset)
);

// actor sub_bytes_5
sub_bytes actor_sub_bytes_5 (
	// Input Signal(s)
	.in_state(sub_bytes_5_in_state_data),
	.in_state_rd(sub_bytes_5_in_state_rd),
	.in_state_empty(sub_bytes_5_in_state_empty)
	,
	
	// Output Signal(s)
	.out_state(sub_bytes_5_out_state_data),
	.out_state_wr(sub_bytes_5_out_state_wr),
	.out_state_full(sub_bytes_5_out_state_full)
		,
	
	// System Signal(s)
	.clock(clock),
	.reset(reset)
);


// fifo_small_shift_rows_5_in_state
fifo_small #(
	.depth(64),
	.size(128)
) fifo_small_shift_rows_5_in_state(
	.datain(fifo_small_shift_rows_5_in_state_data),
	.dataout(shift_rows_5_in_state_data),
	.enr(shift_rows_5_in_state_rd),
	.enw(fifo_small_shift_rows_5_in_state_wr),
	.empty(shift_rows_5_in_state_empty),
	.full(fifo_small_shift_rows_5_in_state_full),
	
	// System Signal(s)
	.clk(clock),
	.rst(reset)
);

// actor shift_rows_5
shift_rows actor_shift_rows_5 (
	// Input Signal(s)
	.in_state(shift_rows_5_in_state_data),
	.in_state_rd(shift_rows_5_in_state_rd),
	.in_state_empty(shift_rows_5_in_state_empty)
	,
	
	// Output Signal(s)
	.out_state(shift_rows_5_out_state_data),
	.out_state_wr(shift_rows_5_out_state_wr),
	.out_state_full(shift_rows_5_out_state_full)
		,
	
	// System Signal(s)
	.clock(clock),
	.reset(reset)
);


// fifo_small_mix_cols_4_in_state
fifo_small #(
	.depth(64),
	.size(128)
) fifo_small_mix_cols_4_in_state(
	.datain(fifo_small_mix_cols_4_in_state_data),
	.dataout(mix_cols_4_in_state_data),
	.enr(mix_cols_4_in_state_rd),
	.enw(fifo_small_mix_cols_4_in_state_wr),
	.empty(mix_cols_4_in_state_empty),
	.full(fifo_small_mix_cols_4_in_state_full),
	
	// System Signal(s)
	.clk(clock),
	.rst(reset)
);

// actor mix_cols_4
mix_cols actor_mix_cols_4 (
	// Input Signal(s)
	.in_state(mix_cols_4_in_state_data),
	.in_state_rd(mix_cols_4_in_state_rd),
	.in_state_empty(mix_cols_4_in_state_empty)
	,
	
	// Output Signal(s)
	.out_state(mix_cols_4_out_state_data),
	.out_state_wr(mix_cols_4_out_state_wr),
	.out_state_full(mix_cols_4_out_state_full)
		,
	
	// System Signal(s)
	.clock(clock),
	.reset(reset)
);


// fifo_small_add_round_key_6_in_state
fifo_small #(
	.depth(64),
	.size(128)
) fifo_small_add_round_key_6_in_state(
	.datain(fifo_small_add_round_key_6_in_state_data),
	.dataout(add_round_key_6_in_state_data),
	.enr(add_round_key_6_in_state_rd),
	.enw(fifo_small_add_round_key_6_in_state_wr),
	.empty(add_round_key_6_in_state_empty),
	.full(fifo_small_add_round_key_6_in_state_full),
	
	// System Signal(s)
	.clk(clock),
	.rst(reset)
);
// fifo_small_add_round_key_6_round_key
fifo_small #(
	.depth(64),
	.size(128)
) fifo_small_add_round_key_6_round_key(
	.datain(fifo_small_add_round_key_6_round_key_data),
	.dataout(add_round_key_6_round_key_data),
	.enr(add_round_key_6_round_key_rd),
	.enw(fifo_small_add_round_key_6_round_key_wr),
	.empty(add_round_key_6_round_key_empty),
	.full(fifo_small_add_round_key_6_round_key_full),
	
	// System Signal(s)
	.clk(clock),
	.rst(reset)
);

// actor add_round_key_6
add_round_key actor_add_round_key_6 (
	// Input Signal(s)
	.in_state(add_round_key_6_in_state_data),
	.in_state_rd(add_round_key_6_in_state_rd),
	.in_state_empty(add_round_key_6_in_state_empty),
	.round_key(add_round_key_6_round_key_data),
	.round_key_rd(add_round_key_6_round_key_rd),
	.round_key_empty(add_round_key_6_round_key_empty)
	,
	
	// Output Signal(s)
	.out_state(add_round_key_6_out_state_data),
	.out_state_wr(add_round_key_6_out_state_wr),
	.out_state_full(add_round_key_6_out_state_full)
		,
	
	// System Signal(s)
	.clock(clock),
	.reset(reset)
);


// fifo_small_sub_bytes_6_in_state
fifo_small #(
	.depth(64),
	.size(128)
) fifo_small_sub_bytes_6_in_state(
	.datain(fifo_small_sub_bytes_6_in_state_data),
	.dataout(sub_bytes_6_in_state_data),
	.enr(sub_bytes_6_in_state_rd),
	.enw(fifo_small_sub_bytes_6_in_state_wr),
	.empty(sub_bytes_6_in_state_empty),
	.full(fifo_small_sub_bytes_6_in_state_full),
	
	// System Signal(s)
	.clk(clock),
	.rst(reset)
);

// actor sub_bytes_6
sub_bytes actor_sub_bytes_6 (
	// Input Signal(s)
	.in_state(sub_bytes_6_in_state_data),
	.in_state_rd(sub_bytes_6_in_state_rd),
	.in_state_empty(sub_bytes_6_in_state_empty)
	,
	
	// Output Signal(s)
	.out_state(sub_bytes_6_out_state_data),
	.out_state_wr(sub_bytes_6_out_state_wr),
	.out_state_full(sub_bytes_6_out_state_full)
		,
	
	// System Signal(s)
	.clock(clock),
	.reset(reset)
);


// fifo_small_shift_rows_6_in_state
fifo_small #(
	.depth(64),
	.size(128)
) fifo_small_shift_rows_6_in_state(
	.datain(fifo_small_shift_rows_6_in_state_data),
	.dataout(shift_rows_6_in_state_data),
	.enr(shift_rows_6_in_state_rd),
	.enw(fifo_small_shift_rows_6_in_state_wr),
	.empty(shift_rows_6_in_state_empty),
	.full(fifo_small_shift_rows_6_in_state_full),
	
	// System Signal(s)
	.clk(clock),
	.rst(reset)
);

// actor shift_rows_6
shift_rows actor_shift_rows_6 (
	// Input Signal(s)
	.in_state(shift_rows_6_in_state_data),
	.in_state_rd(shift_rows_6_in_state_rd),
	.in_state_empty(shift_rows_6_in_state_empty)
	,
	
	// Output Signal(s)
	.out_state(shift_rows_6_out_state_data),
	.out_state_wr(shift_rows_6_out_state_wr),
	.out_state_full(shift_rows_6_out_state_full)
		,
	
	// System Signal(s)
	.clock(clock),
	.reset(reset)
);


// fifo_small_mix_cols_5_in_state
fifo_small #(
	.depth(64),
	.size(128)
) fifo_small_mix_cols_5_in_state(
	.datain(fifo_small_mix_cols_5_in_state_data),
	.dataout(mix_cols_5_in_state_data),
	.enr(mix_cols_5_in_state_rd),
	.enw(fifo_small_mix_cols_5_in_state_wr),
	.empty(mix_cols_5_in_state_empty),
	.full(fifo_small_mix_cols_5_in_state_full),
	
	// System Signal(s)
	.clk(clock),
	.rst(reset)
);

// actor mix_cols_5
mix_cols actor_mix_cols_5 (
	// Input Signal(s)
	.in_state(mix_cols_5_in_state_data),
	.in_state_rd(mix_cols_5_in_state_rd),
	.in_state_empty(mix_cols_5_in_state_empty)
	,
	
	// Output Signal(s)
	.out_state(mix_cols_5_out_state_data),
	.out_state_wr(mix_cols_5_out_state_wr),
	.out_state_full(mix_cols_5_out_state_full)
		,
	
	// System Signal(s)
	.clock(clock),
	.reset(reset)
);


// fifo_small_add_round_key_7_in_state
fifo_small #(
	.depth(64),
	.size(128)
) fifo_small_add_round_key_7_in_state(
	.datain(fifo_small_add_round_key_7_in_state_data),
	.dataout(add_round_key_7_in_state_data),
	.enr(add_round_key_7_in_state_rd),
	.enw(fifo_small_add_round_key_7_in_state_wr),
	.empty(add_round_key_7_in_state_empty),
	.full(fifo_small_add_round_key_7_in_state_full),
	
	// System Signal(s)
	.clk(clock),
	.rst(reset)
);
// fifo_small_add_round_key_7_round_key
fifo_small #(
	.depth(64),
	.size(128)
) fifo_small_add_round_key_7_round_key(
	.datain(fifo_small_add_round_key_7_round_key_data),
	.dataout(add_round_key_7_round_key_data),
	.enr(add_round_key_7_round_key_rd),
	.enw(fifo_small_add_round_key_7_round_key_wr),
	.empty(add_round_key_7_round_key_empty),
	.full(fifo_small_add_round_key_7_round_key_full),
	
	// System Signal(s)
	.clk(clock),
	.rst(reset)
);

// actor add_round_key_7
add_round_key actor_add_round_key_7 (
	// Input Signal(s)
	.in_state(add_round_key_7_in_state_data),
	.in_state_rd(add_round_key_7_in_state_rd),
	.in_state_empty(add_round_key_7_in_state_empty),
	.round_key(add_round_key_7_round_key_data),
	.round_key_rd(add_round_key_7_round_key_rd),
	.round_key_empty(add_round_key_7_round_key_empty)
	,
	
	// Output Signal(s)
	.out_state(add_round_key_7_out_state_data),
	.out_state_wr(add_round_key_7_out_state_wr),
	.out_state_full(add_round_key_7_out_state_full)
		,
	
	// System Signal(s)
	.clock(clock),
	.reset(reset)
);


// fifo_small_sub_bytes_7_in_state
fifo_small #(
	.depth(64),
	.size(128)
) fifo_small_sub_bytes_7_in_state(
	.datain(fifo_small_sub_bytes_7_in_state_data),
	.dataout(sub_bytes_7_in_state_data),
	.enr(sub_bytes_7_in_state_rd),
	.enw(fifo_small_sub_bytes_7_in_state_wr),
	.empty(sub_bytes_7_in_state_empty),
	.full(fifo_small_sub_bytes_7_in_state_full),
	
	// System Signal(s)
	.clk(clock),
	.rst(reset)
);

// actor sub_bytes_7
sub_bytes actor_sub_bytes_7 (
	// Input Signal(s)
	.in_state(sub_bytes_7_in_state_data),
	.in_state_rd(sub_bytes_7_in_state_rd),
	.in_state_empty(sub_bytes_7_in_state_empty)
	,
	
	// Output Signal(s)
	.out_state(sub_bytes_7_out_state_data),
	.out_state_wr(sub_bytes_7_out_state_wr),
	.out_state_full(sub_bytes_7_out_state_full)
		,
	
	// System Signal(s)
	.clock(clock),
	.reset(reset)
);


// fifo_small_shift_rows_7_in_state
fifo_small #(
	.depth(64),
	.size(128)
) fifo_small_shift_rows_7_in_state(
	.datain(fifo_small_shift_rows_7_in_state_data),
	.dataout(shift_rows_7_in_state_data),
	.enr(shift_rows_7_in_state_rd),
	.enw(fifo_small_shift_rows_7_in_state_wr),
	.empty(shift_rows_7_in_state_empty),
	.full(fifo_small_shift_rows_7_in_state_full),
	
	// System Signal(s)
	.clk(clock),
	.rst(reset)
);

// actor shift_rows_7
shift_rows actor_shift_rows_7 (
	// Input Signal(s)
	.in_state(shift_rows_7_in_state_data),
	.in_state_rd(shift_rows_7_in_state_rd),
	.in_state_empty(shift_rows_7_in_state_empty)
	,
	
	// Output Signal(s)
	.out_state(shift_rows_7_out_state_data),
	.out_state_wr(shift_rows_7_out_state_wr),
	.out_state_full(shift_rows_7_out_state_full)
		,
	
	// System Signal(s)
	.clock(clock),
	.reset(reset)
);


// fifo_small_mix_cols_6_in_state
fifo_small #(
	.depth(64),
	.size(128)
) fifo_small_mix_cols_6_in_state(
	.datain(fifo_small_mix_cols_6_in_state_data),
	.dataout(mix_cols_6_in_state_data),
	.enr(mix_cols_6_in_state_rd),
	.enw(fifo_small_mix_cols_6_in_state_wr),
	.empty(mix_cols_6_in_state_empty),
	.full(fifo_small_mix_cols_6_in_state_full),
	
	// System Signal(s)
	.clk(clock),
	.rst(reset)
);

// actor mix_cols_6
mix_cols actor_mix_cols_6 (
	// Input Signal(s)
	.in_state(mix_cols_6_in_state_data),
	.in_state_rd(mix_cols_6_in_state_rd),
	.in_state_empty(mix_cols_6_in_state_empty)
	,
	
	// Output Signal(s)
	.out_state(mix_cols_6_out_state_data),
	.out_state_wr(mix_cols_6_out_state_wr),
	.out_state_full(mix_cols_6_out_state_full)
		,
	
	// System Signal(s)
	.clock(clock),
	.reset(reset)
);


// fifo_small_add_round_key_8_in_state
fifo_small #(
	.depth(64),
	.size(128)
) fifo_small_add_round_key_8_in_state(
	.datain(fifo_small_add_round_key_8_in_state_data),
	.dataout(add_round_key_8_in_state_data),
	.enr(add_round_key_8_in_state_rd),
	.enw(fifo_small_add_round_key_8_in_state_wr),
	.empty(add_round_key_8_in_state_empty),
	.full(fifo_small_add_round_key_8_in_state_full),
	
	// System Signal(s)
	.clk(clock),
	.rst(reset)
);
// fifo_small_add_round_key_8_round_key
fifo_small #(
	.depth(64),
	.size(128)
) fifo_small_add_round_key_8_round_key(
	.datain(fifo_small_add_round_key_8_round_key_data),
	.dataout(add_round_key_8_round_key_data),
	.enr(add_round_key_8_round_key_rd),
	.enw(fifo_small_add_round_key_8_round_key_wr),
	.empty(add_round_key_8_round_key_empty),
	.full(fifo_small_add_round_key_8_round_key_full),
	
	// System Signal(s)
	.clk(clock),
	.rst(reset)
);

// actor add_round_key_8
add_round_key actor_add_round_key_8 (
	// Input Signal(s)
	.in_state(add_round_key_8_in_state_data),
	.in_state_rd(add_round_key_8_in_state_rd),
	.in_state_empty(add_round_key_8_in_state_empty),
	.round_key(add_round_key_8_round_key_data),
	.round_key_rd(add_round_key_8_round_key_rd),
	.round_key_empty(add_round_key_8_round_key_empty)
	,
	
	// Output Signal(s)
	.out_state(add_round_key_8_out_state_data),
	.out_state_wr(add_round_key_8_out_state_wr),
	.out_state_full(add_round_key_8_out_state_full)
		,
	
	// System Signal(s)
	.clock(clock),
	.reset(reset)
);


// fifo_small_sub_bytes_8_in_state
fifo_small #(
	.depth(64),
	.size(128)
) fifo_small_sub_bytes_8_in_state(
	.datain(fifo_small_sub_bytes_8_in_state_data),
	.dataout(sub_bytes_8_in_state_data),
	.enr(sub_bytes_8_in_state_rd),
	.enw(fifo_small_sub_bytes_8_in_state_wr),
	.empty(sub_bytes_8_in_state_empty),
	.full(fifo_small_sub_bytes_8_in_state_full),
	
	// System Signal(s)
	.clk(clock),
	.rst(reset)
);

// actor sub_bytes_8
sub_bytes actor_sub_bytes_8 (
	// Input Signal(s)
	.in_state(sub_bytes_8_in_state_data),
	.in_state_rd(sub_bytes_8_in_state_rd),
	.in_state_empty(sub_bytes_8_in_state_empty)
	,
	
	// Output Signal(s)
	.out_state(sub_bytes_8_out_state_data),
	.out_state_wr(sub_bytes_8_out_state_wr),
	.out_state_full(sub_bytes_8_out_state_full)
		,
	
	// System Signal(s)
	.clock(clock),
	.reset(reset)
);


// fifo_small_shift_rows_8_in_state
fifo_small #(
	.depth(64),
	.size(128)
) fifo_small_shift_rows_8_in_state(
	.datain(fifo_small_shift_rows_8_in_state_data),
	.dataout(shift_rows_8_in_state_data),
	.enr(shift_rows_8_in_state_rd),
	.enw(fifo_small_shift_rows_8_in_state_wr),
	.empty(shift_rows_8_in_state_empty),
	.full(fifo_small_shift_rows_8_in_state_full),
	
	// System Signal(s)
	.clk(clock),
	.rst(reset)
);

// actor shift_rows_8
shift_rows actor_shift_rows_8 (
	// Input Signal(s)
	.in_state(shift_rows_8_in_state_data),
	.in_state_rd(shift_rows_8_in_state_rd),
	.in_state_empty(shift_rows_8_in_state_empty)
	,
	
	// Output Signal(s)
	.out_state(shift_rows_8_out_state_data),
	.out_state_wr(shift_rows_8_out_state_wr),
	.out_state_full(shift_rows_8_out_state_full)
		,
	
	// System Signal(s)
	.clock(clock),
	.reset(reset)
);


// fifo_small_mix_cols_7_in_state
fifo_small #(
	.depth(64),
	.size(128)
) fifo_small_mix_cols_7_in_state(
	.datain(fifo_small_mix_cols_7_in_state_data),
	.dataout(mix_cols_7_in_state_data),
	.enr(mix_cols_7_in_state_rd),
	.enw(fifo_small_mix_cols_7_in_state_wr),
	.empty(mix_cols_7_in_state_empty),
	.full(fifo_small_mix_cols_7_in_state_full),
	
	// System Signal(s)
	.clk(clock),
	.rst(reset)
);

// actor mix_cols_7
mix_cols actor_mix_cols_7 (
	// Input Signal(s)
	.in_state(mix_cols_7_in_state_data),
	.in_state_rd(mix_cols_7_in_state_rd),
	.in_state_empty(mix_cols_7_in_state_empty)
	,
	
	// Output Signal(s)
	.out_state(mix_cols_7_out_state_data),
	.out_state_wr(mix_cols_7_out_state_wr),
	.out_state_full(mix_cols_7_out_state_full)
		,
	
	// System Signal(s)
	.clock(clock),
	.reset(reset)
);


// fifo_small_add_round_key_9_in_state
fifo_small #(
	.depth(64),
	.size(128)
) fifo_small_add_round_key_9_in_state(
	.datain(fifo_small_add_round_key_9_in_state_data),
	.dataout(add_round_key_9_in_state_data),
	.enr(add_round_key_9_in_state_rd),
	.enw(fifo_small_add_round_key_9_in_state_wr),
	.empty(add_round_key_9_in_state_empty),
	.full(fifo_small_add_round_key_9_in_state_full),
	
	// System Signal(s)
	.clk(clock),
	.rst(reset)
);
// fifo_small_add_round_key_9_round_key
fifo_small #(
	.depth(64),
	.size(128)
) fifo_small_add_round_key_9_round_key(
	.datain(fifo_small_add_round_key_9_round_key_data),
	.dataout(add_round_key_9_round_key_data),
	.enr(add_round_key_9_round_key_rd),
	.enw(fifo_small_add_round_key_9_round_key_wr),
	.empty(add_round_key_9_round_key_empty),
	.full(fifo_small_add_round_key_9_round_key_full),
	
	// System Signal(s)
	.clk(clock),
	.rst(reset)
);

// actor add_round_key_9
add_round_key actor_add_round_key_9 (
	// Input Signal(s)
	.in_state(add_round_key_9_in_state_data),
	.in_state_rd(add_round_key_9_in_state_rd),
	.in_state_empty(add_round_key_9_in_state_empty),
	.round_key(add_round_key_9_round_key_data),
	.round_key_rd(add_round_key_9_round_key_rd),
	.round_key_empty(add_round_key_9_round_key_empty)
	,
	
	// Output Signal(s)
	.out_state(add_round_key_9_out_state_data),
	.out_state_wr(add_round_key_9_out_state_wr),
	.out_state_full(add_round_key_9_out_state_full)
		,
	
	// System Signal(s)
	.clock(clock),
	.reset(reset)
);


// fifo_small_expand_key0_128_0_in_key
fifo_small #(
	.depth(64),
	.size(128)
) fifo_small_expand_key0_128_0_in_key(
	.datain(fifo_small_expand_key0_128_0_in_key_data),
	.dataout(expand_key0_128_0_in_key_data),
	.enr(expand_key0_128_0_in_key_rd),
	.enw(fifo_small_expand_key0_128_0_in_key_wr),
	.empty(expand_key0_128_0_in_key_empty),
	.full(fifo_small_expand_key0_128_0_in_key_full),
	
	// System Signal(s)
	.clk(clock),
	.rst(reset)
);
// fifo_small_expand_key0_128_0_in_rc
fifo_small #(
	.depth(64),
	.size(8)
) fifo_small_expand_key0_128_0_in_rc(
	.datain(fifo_small_expand_key0_128_0_in_rc_data),
	.dataout(expand_key0_128_0_in_rc_data),
	.enr(expand_key0_128_0_in_rc_rd),
	.enw(fifo_small_expand_key0_128_0_in_rc_wr),
	.empty(expand_key0_128_0_in_rc_empty),
	.full(fifo_small_expand_key0_128_0_in_rc_full),
	
	// System Signal(s)
	.clk(clock),
	.rst(reset)
);

// actor expand_key0_128_0
expand_key0_128 actor_expand_key0_128_0 (
	// Input Signal(s)
	.in_key(expand_key0_128_0_in_key_data),
	.in_key_rd(expand_key0_128_0_in_key_rd),
	.in_key_empty(expand_key0_128_0_in_key_empty),
	.in_rc(expand_key0_128_0_in_rc_data),
	.in_rc_rd(expand_key0_128_0_in_rc_rd),
	.in_rc_empty(expand_key0_128_0_in_rc_empty)
	,
	
	// Output Signal(s)
	.out_key(expand_key0_128_0_out_key_data),
	.out_key_wr(expand_key0_128_0_out_key_wr),
	.out_key_full(expand_key0_128_0_out_key_full)
		,
	
	// System Signal(s)
	.clock(clock),
	.reset(reset)
);


// fifo_small_expand_key1_128_0_in_key
fifo_small #(
	.depth(64),
	.size(128)
) fifo_small_expand_key1_128_0_in_key(
	.datain(fifo_small_expand_key1_128_0_in_key_data),
	.dataout(expand_key1_128_0_in_key_data),
	.enr(expand_key1_128_0_in_key_rd),
	.enw(fifo_small_expand_key1_128_0_in_key_wr),
	.empty(expand_key1_128_0_in_key_empty),
	.full(fifo_small_expand_key1_128_0_in_key_full),
	
	// System Signal(s)
	.clk(clock),
	.rst(reset)
);

// actor expand_key1_128_0
expand_key1_128 actor_expand_key1_128_0 (
	// Input Signal(s)
	.in_key(expand_key1_128_0_in_key_data),
	.in_key_rd(expand_key1_128_0_in_key_rd),
	.in_key_empty(expand_key1_128_0_in_key_empty)
	,
	
	// Output Signal(s)
	.out_key(expand_key1_128_0_out_key_data),
	.out_key_wr(expand_key1_128_0_out_key_wr),
	.out_key_full(expand_key1_128_0_out_key_full)
		,
	
	// System Signal(s)
	.clock(clock),
	.reset(reset)
);


// fifo_small_expand_key2_128_0_in_key
fifo_small #(
	.depth(64),
	.size(128)
) fifo_small_expand_key2_128_0_in_key(
	.datain(fifo_small_expand_key2_128_0_in_key_data),
	.dataout(expand_key2_128_0_in_key_data),
	.enr(expand_key2_128_0_in_key_rd),
	.enw(fifo_small_expand_key2_128_0_in_key_wr),
	.empty(expand_key2_128_0_in_key_empty),
	.full(fifo_small_expand_key2_128_0_in_key_full),
	
	// System Signal(s)
	.clk(clock),
	.rst(reset)
);

// actor expand_key2_128_0
expand_key2_128 actor_expand_key2_128_0 (
	// Input Signal(s)
	.in_key(expand_key2_128_0_in_key_data),
	.in_key_rd(expand_key2_128_0_in_key_rd),
	.in_key_empty(expand_key2_128_0_in_key_empty)
	,
	
	// Output Signal(s)
	.out_key(expand_key2_128_0_out_key_data),
	.out_key_wr(expand_key2_128_0_out_key_wr),
	.out_key_full(expand_key2_128_0_out_key_full)
		,
	
	// System Signal(s)
	.clock(clock),
	.reset(reset)
);


// fifo_small_expand_key3_128_0_in_key
fifo_small #(
	.depth(64),
	.size(128)
) fifo_small_expand_key3_128_0_in_key(
	.datain(fifo_small_expand_key3_128_0_in_key_data),
	.dataout(expand_key3_128_0_in_key_data),
	.enr(expand_key3_128_0_in_key_rd),
	.enw(fifo_small_expand_key3_128_0_in_key_wr),
	.empty(expand_key3_128_0_in_key_empty),
	.full(fifo_small_expand_key3_128_0_in_key_full),
	
	// System Signal(s)
	.clk(clock),
	.rst(reset)
);

// actor expand_key3_128_0
expand_key3_128 actor_expand_key3_128_0 (
	// Input Signal(s)
	.in_key(expand_key3_128_0_in_key_data),
	.in_key_rd(expand_key3_128_0_in_key_rd),
	.in_key_empty(expand_key3_128_0_in_key_empty)
	,
	
	// Output Signal(s)
	.out_key(expand_key3_128_0_out_key_data),
	.out_key_wr(expand_key3_128_0_out_key_wr),
	.out_key_full(expand_key3_128_0_out_key_full)
		,
	
	// System Signal(s)
	.clock(clock),
	.reset(reset)
);


// fifo_small_expand_key0_128_1_in_key
fifo_small #(
	.depth(64),
	.size(128)
) fifo_small_expand_key0_128_1_in_key(
	.datain(fifo_small_expand_key0_128_1_in_key_data),
	.dataout(expand_key0_128_1_in_key_data),
	.enr(expand_key0_128_1_in_key_rd),
	.enw(fifo_small_expand_key0_128_1_in_key_wr),
	.empty(expand_key0_128_1_in_key_empty),
	.full(fifo_small_expand_key0_128_1_in_key_full),
	
	// System Signal(s)
	.clk(clock),
	.rst(reset)
);
// fifo_small_expand_key0_128_1_in_rc
fifo_small #(
	.depth(64),
	.size(8)
) fifo_small_expand_key0_128_1_in_rc(
	.datain(fifo_small_expand_key0_128_1_in_rc_data),
	.dataout(expand_key0_128_1_in_rc_data),
	.enr(expand_key0_128_1_in_rc_rd),
	.enw(fifo_small_expand_key0_128_1_in_rc_wr),
	.empty(expand_key0_128_1_in_rc_empty),
	.full(fifo_small_expand_key0_128_1_in_rc_full),
	
	// System Signal(s)
	.clk(clock),
	.rst(reset)
);

// actor expand_key0_128_1
expand_key0_128 actor_expand_key0_128_1 (
	// Input Signal(s)
	.in_key(expand_key0_128_1_in_key_data),
	.in_key_rd(expand_key0_128_1_in_key_rd),
	.in_key_empty(expand_key0_128_1_in_key_empty),
	.in_rc(expand_key0_128_1_in_rc_data),
	.in_rc_rd(expand_key0_128_1_in_rc_rd),
	.in_rc_empty(expand_key0_128_1_in_rc_empty)
	,
	
	// Output Signal(s)
	.out_key(expand_key0_128_1_out_key_data),
	.out_key_wr(expand_key0_128_1_out_key_wr),
	.out_key_full(expand_key0_128_1_out_key_full)
		,
	
	// System Signal(s)
	.clock(clock),
	.reset(reset)
);


// fifo_small_expand_key1_128_1_in_key
fifo_small #(
	.depth(64),
	.size(128)
) fifo_small_expand_key1_128_1_in_key(
	.datain(fifo_small_expand_key1_128_1_in_key_data),
	.dataout(expand_key1_128_1_in_key_data),
	.enr(expand_key1_128_1_in_key_rd),
	.enw(fifo_small_expand_key1_128_1_in_key_wr),
	.empty(expand_key1_128_1_in_key_empty),
	.full(fifo_small_expand_key1_128_1_in_key_full),
	
	// System Signal(s)
	.clk(clock),
	.rst(reset)
);

// actor expand_key1_128_1
expand_key1_128 actor_expand_key1_128_1 (
	// Input Signal(s)
	.in_key(expand_key1_128_1_in_key_data),
	.in_key_rd(expand_key1_128_1_in_key_rd),
	.in_key_empty(expand_key1_128_1_in_key_empty)
	,
	
	// Output Signal(s)
	.out_key(expand_key1_128_1_out_key_data),
	.out_key_wr(expand_key1_128_1_out_key_wr),
	.out_key_full(expand_key1_128_1_out_key_full)
		,
	
	// System Signal(s)
	.clock(clock),
	.reset(reset)
);


// fifo_small_expand_key2_128_1_in_key
fifo_small #(
	.depth(64),
	.size(128)
) fifo_small_expand_key2_128_1_in_key(
	.datain(fifo_small_expand_key2_128_1_in_key_data),
	.dataout(expand_key2_128_1_in_key_data),
	.enr(expand_key2_128_1_in_key_rd),
	.enw(fifo_small_expand_key2_128_1_in_key_wr),
	.empty(expand_key2_128_1_in_key_empty),
	.full(fifo_small_expand_key2_128_1_in_key_full),
	
	// System Signal(s)
	.clk(clock),
	.rst(reset)
);

// actor expand_key2_128_1
expand_key2_128 actor_expand_key2_128_1 (
	// Input Signal(s)
	.in_key(expand_key2_128_1_in_key_data),
	.in_key_rd(expand_key2_128_1_in_key_rd),
	.in_key_empty(expand_key2_128_1_in_key_empty)
	,
	
	// Output Signal(s)
	.out_key(expand_key2_128_1_out_key_data),
	.out_key_wr(expand_key2_128_1_out_key_wr),
	.out_key_full(expand_key2_128_1_out_key_full)
		,
	
	// System Signal(s)
	.clock(clock),
	.reset(reset)
);


// fifo_small_expand_key3_128_1_in_key
fifo_small #(
	.depth(64),
	.size(128)
) fifo_small_expand_key3_128_1_in_key(
	.datain(fifo_small_expand_key3_128_1_in_key_data),
	.dataout(expand_key3_128_1_in_key_data),
	.enr(expand_key3_128_1_in_key_rd),
	.enw(fifo_small_expand_key3_128_1_in_key_wr),
	.empty(expand_key3_128_1_in_key_empty),
	.full(fifo_small_expand_key3_128_1_in_key_full),
	
	// System Signal(s)
	.clk(clock),
	.rst(reset)
);

// actor expand_key3_128_1
expand_key3_128 actor_expand_key3_128_1 (
	// Input Signal(s)
	.in_key(expand_key3_128_1_in_key_data),
	.in_key_rd(expand_key3_128_1_in_key_rd),
	.in_key_empty(expand_key3_128_1_in_key_empty)
	,
	
	// Output Signal(s)
	.out_key(expand_key3_128_1_out_key_data),
	.out_key_wr(expand_key3_128_1_out_key_wr),
	.out_key_full(expand_key3_128_1_out_key_full)
		,
	
	// System Signal(s)
	.clock(clock),
	.reset(reset)
);


// fifo_small_expand_key0_128_2_in_key
fifo_small #(
	.depth(64),
	.size(128)
) fifo_small_expand_key0_128_2_in_key(
	.datain(fifo_small_expand_key0_128_2_in_key_data),
	.dataout(expand_key0_128_2_in_key_data),
	.enr(expand_key0_128_2_in_key_rd),
	.enw(fifo_small_expand_key0_128_2_in_key_wr),
	.empty(expand_key0_128_2_in_key_empty),
	.full(fifo_small_expand_key0_128_2_in_key_full),
	
	// System Signal(s)
	.clk(clock),
	.rst(reset)
);
// fifo_small_expand_key0_128_2_in_rc
fifo_small #(
	.depth(64),
	.size(8)
) fifo_small_expand_key0_128_2_in_rc(
	.datain(fifo_small_expand_key0_128_2_in_rc_data),
	.dataout(expand_key0_128_2_in_rc_data),
	.enr(expand_key0_128_2_in_rc_rd),
	.enw(fifo_small_expand_key0_128_2_in_rc_wr),
	.empty(expand_key0_128_2_in_rc_empty),
	.full(fifo_small_expand_key0_128_2_in_rc_full),
	
	// System Signal(s)
	.clk(clock),
	.rst(reset)
);

// actor expand_key0_128_2
expand_key0_128 actor_expand_key0_128_2 (
	// Input Signal(s)
	.in_key(expand_key0_128_2_in_key_data),
	.in_key_rd(expand_key0_128_2_in_key_rd),
	.in_key_empty(expand_key0_128_2_in_key_empty),
	.in_rc(expand_key0_128_2_in_rc_data),
	.in_rc_rd(expand_key0_128_2_in_rc_rd),
	.in_rc_empty(expand_key0_128_2_in_rc_empty)
	,
	
	// Output Signal(s)
	.out_key(expand_key0_128_2_out_key_data),
	.out_key_wr(expand_key0_128_2_out_key_wr),
	.out_key_full(expand_key0_128_2_out_key_full)
		,
	
	// System Signal(s)
	.clock(clock),
	.reset(reset)
);


// fifo_small_expand_key1_128_2_in_key
fifo_small #(
	.depth(64),
	.size(128)
) fifo_small_expand_key1_128_2_in_key(
	.datain(fifo_small_expand_key1_128_2_in_key_data),
	.dataout(expand_key1_128_2_in_key_data),
	.enr(expand_key1_128_2_in_key_rd),
	.enw(fifo_small_expand_key1_128_2_in_key_wr),
	.empty(expand_key1_128_2_in_key_empty),
	.full(fifo_small_expand_key1_128_2_in_key_full),
	
	// System Signal(s)
	.clk(clock),
	.rst(reset)
);

// actor expand_key1_128_2
expand_key1_128 actor_expand_key1_128_2 (
	// Input Signal(s)
	.in_key(expand_key1_128_2_in_key_data),
	.in_key_rd(expand_key1_128_2_in_key_rd),
	.in_key_empty(expand_key1_128_2_in_key_empty)
	,
	
	// Output Signal(s)
	.out_key(expand_key1_128_2_out_key_data),
	.out_key_wr(expand_key1_128_2_out_key_wr),
	.out_key_full(expand_key1_128_2_out_key_full)
		,
	
	// System Signal(s)
	.clock(clock),
	.reset(reset)
);


// fifo_small_expand_key2_128_2_in_key
fifo_small #(
	.depth(64),
	.size(128)
) fifo_small_expand_key2_128_2_in_key(
	.datain(fifo_small_expand_key2_128_2_in_key_data),
	.dataout(expand_key2_128_2_in_key_data),
	.enr(expand_key2_128_2_in_key_rd),
	.enw(fifo_small_expand_key2_128_2_in_key_wr),
	.empty(expand_key2_128_2_in_key_empty),
	.full(fifo_small_expand_key2_128_2_in_key_full),
	
	// System Signal(s)
	.clk(clock),
	.rst(reset)
);

// actor expand_key2_128_2
expand_key2_128 actor_expand_key2_128_2 (
	// Input Signal(s)
	.in_key(expand_key2_128_2_in_key_data),
	.in_key_rd(expand_key2_128_2_in_key_rd),
	.in_key_empty(expand_key2_128_2_in_key_empty)
	,
	
	// Output Signal(s)
	.out_key(expand_key2_128_2_out_key_data),
	.out_key_wr(expand_key2_128_2_out_key_wr),
	.out_key_full(expand_key2_128_2_out_key_full)
		,
	
	// System Signal(s)
	.clock(clock),
	.reset(reset)
);


// fifo_small_expand_key3_128_2_in_key
fifo_small #(
	.depth(64),
	.size(128)
) fifo_small_expand_key3_128_2_in_key(
	.datain(fifo_small_expand_key3_128_2_in_key_data),
	.dataout(expand_key3_128_2_in_key_data),
	.enr(expand_key3_128_2_in_key_rd),
	.enw(fifo_small_expand_key3_128_2_in_key_wr),
	.empty(expand_key3_128_2_in_key_empty),
	.full(fifo_small_expand_key3_128_2_in_key_full),
	
	// System Signal(s)
	.clk(clock),
	.rst(reset)
);

// actor expand_key3_128_2
expand_key3_128 actor_expand_key3_128_2 (
	// Input Signal(s)
	.in_key(expand_key3_128_2_in_key_data),
	.in_key_rd(expand_key3_128_2_in_key_rd),
	.in_key_empty(expand_key3_128_2_in_key_empty)
	,
	
	// Output Signal(s)
	.out_key(expand_key3_128_2_out_key_data),
	.out_key_wr(expand_key3_128_2_out_key_wr),
	.out_key_full(expand_key3_128_2_out_key_full)
		,
	
	// System Signal(s)
	.clock(clock),
	.reset(reset)
);


// fifo_small_expand_key0_128_3_in_key
fifo_small #(
	.depth(64),
	.size(128)
) fifo_small_expand_key0_128_3_in_key(
	.datain(fifo_small_expand_key0_128_3_in_key_data),
	.dataout(expand_key0_128_3_in_key_data),
	.enr(expand_key0_128_3_in_key_rd),
	.enw(fifo_small_expand_key0_128_3_in_key_wr),
	.empty(expand_key0_128_3_in_key_empty),
	.full(fifo_small_expand_key0_128_3_in_key_full),
	
	// System Signal(s)
	.clk(clock),
	.rst(reset)
);
// fifo_small_expand_key0_128_3_in_rc
fifo_small #(
	.depth(64),
	.size(8)
) fifo_small_expand_key0_128_3_in_rc(
	.datain(fifo_small_expand_key0_128_3_in_rc_data),
	.dataout(expand_key0_128_3_in_rc_data),
	.enr(expand_key0_128_3_in_rc_rd),
	.enw(fifo_small_expand_key0_128_3_in_rc_wr),
	.empty(expand_key0_128_3_in_rc_empty),
	.full(fifo_small_expand_key0_128_3_in_rc_full),
	
	// System Signal(s)
	.clk(clock),
	.rst(reset)
);

// actor expand_key0_128_3
expand_key0_128 actor_expand_key0_128_3 (
	// Input Signal(s)
	.in_key(expand_key0_128_3_in_key_data),
	.in_key_rd(expand_key0_128_3_in_key_rd),
	.in_key_empty(expand_key0_128_3_in_key_empty),
	.in_rc(expand_key0_128_3_in_rc_data),
	.in_rc_rd(expand_key0_128_3_in_rc_rd),
	.in_rc_empty(expand_key0_128_3_in_rc_empty)
	,
	
	// Output Signal(s)
	.out_key(expand_key0_128_3_out_key_data),
	.out_key_wr(expand_key0_128_3_out_key_wr),
	.out_key_full(expand_key0_128_3_out_key_full)
		,
	
	// System Signal(s)
	.clock(clock),
	.reset(reset)
);


// fifo_small_expand_key1_128_3_in_key
fifo_small #(
	.depth(64),
	.size(128)
) fifo_small_expand_key1_128_3_in_key(
	.datain(fifo_small_expand_key1_128_3_in_key_data),
	.dataout(expand_key1_128_3_in_key_data),
	.enr(expand_key1_128_3_in_key_rd),
	.enw(fifo_small_expand_key1_128_3_in_key_wr),
	.empty(expand_key1_128_3_in_key_empty),
	.full(fifo_small_expand_key1_128_3_in_key_full),
	
	// System Signal(s)
	.clk(clock),
	.rst(reset)
);

// actor expand_key1_128_3
expand_key1_128 actor_expand_key1_128_3 (
	// Input Signal(s)
	.in_key(expand_key1_128_3_in_key_data),
	.in_key_rd(expand_key1_128_3_in_key_rd),
	.in_key_empty(expand_key1_128_3_in_key_empty)
	,
	
	// Output Signal(s)
	.out_key(expand_key1_128_3_out_key_data),
	.out_key_wr(expand_key1_128_3_out_key_wr),
	.out_key_full(expand_key1_128_3_out_key_full)
		,
	
	// System Signal(s)
	.clock(clock),
	.reset(reset)
);


// fifo_small_expand_key2_128_3_in_key
fifo_small #(
	.depth(64),
	.size(128)
) fifo_small_expand_key2_128_3_in_key(
	.datain(fifo_small_expand_key2_128_3_in_key_data),
	.dataout(expand_key2_128_3_in_key_data),
	.enr(expand_key2_128_3_in_key_rd),
	.enw(fifo_small_expand_key2_128_3_in_key_wr),
	.empty(expand_key2_128_3_in_key_empty),
	.full(fifo_small_expand_key2_128_3_in_key_full),
	
	// System Signal(s)
	.clk(clock),
	.rst(reset)
);

// actor expand_key2_128_3
expand_key2_128 actor_expand_key2_128_3 (
	// Input Signal(s)
	.in_key(expand_key2_128_3_in_key_data),
	.in_key_rd(expand_key2_128_3_in_key_rd),
	.in_key_empty(expand_key2_128_3_in_key_empty)
	,
	
	// Output Signal(s)
	.out_key(expand_key2_128_3_out_key_data),
	.out_key_wr(expand_key2_128_3_out_key_wr),
	.out_key_full(expand_key2_128_3_out_key_full)
		,
	
	// System Signal(s)
	.clock(clock),
	.reset(reset)
);


// fifo_small_expand_key3_128_3_in_key
fifo_small #(
	.depth(64),
	.size(128)
) fifo_small_expand_key3_128_3_in_key(
	.datain(fifo_small_expand_key3_128_3_in_key_data),
	.dataout(expand_key3_128_3_in_key_data),
	.enr(expand_key3_128_3_in_key_rd),
	.enw(fifo_small_expand_key3_128_3_in_key_wr),
	.empty(expand_key3_128_3_in_key_empty),
	.full(fifo_small_expand_key3_128_3_in_key_full),
	
	// System Signal(s)
	.clk(clock),
	.rst(reset)
);

// actor expand_key3_128_3
expand_key3_128 actor_expand_key3_128_3 (
	// Input Signal(s)
	.in_key(expand_key3_128_3_in_key_data),
	.in_key_rd(expand_key3_128_3_in_key_rd),
	.in_key_empty(expand_key3_128_3_in_key_empty)
	,
	
	// Output Signal(s)
	.out_key(expand_key3_128_3_out_key_data),
	.out_key_wr(expand_key3_128_3_out_key_wr),
	.out_key_full(expand_key3_128_3_out_key_full)
		,
	
	// System Signal(s)
	.clock(clock),
	.reset(reset)
);


// fifo_small_expand_key0_128_4_in_key
fifo_small #(
	.depth(64),
	.size(128)
) fifo_small_expand_key0_128_4_in_key(
	.datain(fifo_small_expand_key0_128_4_in_key_data),
	.dataout(expand_key0_128_4_in_key_data),
	.enr(expand_key0_128_4_in_key_rd),
	.enw(fifo_small_expand_key0_128_4_in_key_wr),
	.empty(expand_key0_128_4_in_key_empty),
	.full(fifo_small_expand_key0_128_4_in_key_full),
	
	// System Signal(s)
	.clk(clock),
	.rst(reset)
);
// fifo_small_expand_key0_128_4_in_rc
fifo_small #(
	.depth(64),
	.size(8)
) fifo_small_expand_key0_128_4_in_rc(
	.datain(fifo_small_expand_key0_128_4_in_rc_data),
	.dataout(expand_key0_128_4_in_rc_data),
	.enr(expand_key0_128_4_in_rc_rd),
	.enw(fifo_small_expand_key0_128_4_in_rc_wr),
	.empty(expand_key0_128_4_in_rc_empty),
	.full(fifo_small_expand_key0_128_4_in_rc_full),
	
	// System Signal(s)
	.clk(clock),
	.rst(reset)
);

// actor expand_key0_128_4
expand_key0_128 actor_expand_key0_128_4 (
	// Input Signal(s)
	.in_key(expand_key0_128_4_in_key_data),
	.in_key_rd(expand_key0_128_4_in_key_rd),
	.in_key_empty(expand_key0_128_4_in_key_empty),
	.in_rc(expand_key0_128_4_in_rc_data),
	.in_rc_rd(expand_key0_128_4_in_rc_rd),
	.in_rc_empty(expand_key0_128_4_in_rc_empty)
	,
	
	// Output Signal(s)
	.out_key(expand_key0_128_4_out_key_data),
	.out_key_wr(expand_key0_128_4_out_key_wr),
	.out_key_full(expand_key0_128_4_out_key_full)
		,
	
	// System Signal(s)
	.clock(clock),
	.reset(reset)
);


// fifo_small_expand_key1_128_4_in_key
fifo_small #(
	.depth(64),
	.size(128)
) fifo_small_expand_key1_128_4_in_key(
	.datain(fifo_small_expand_key1_128_4_in_key_data),
	.dataout(expand_key1_128_4_in_key_data),
	.enr(expand_key1_128_4_in_key_rd),
	.enw(fifo_small_expand_key1_128_4_in_key_wr),
	.empty(expand_key1_128_4_in_key_empty),
	.full(fifo_small_expand_key1_128_4_in_key_full),
	
	// System Signal(s)
	.clk(clock),
	.rst(reset)
);

// actor expand_key1_128_4
expand_key1_128 actor_expand_key1_128_4 (
	// Input Signal(s)
	.in_key(expand_key1_128_4_in_key_data),
	.in_key_rd(expand_key1_128_4_in_key_rd),
	.in_key_empty(expand_key1_128_4_in_key_empty)
	,
	
	// Output Signal(s)
	.out_key(expand_key1_128_4_out_key_data),
	.out_key_wr(expand_key1_128_4_out_key_wr),
	.out_key_full(expand_key1_128_4_out_key_full)
		,
	
	// System Signal(s)
	.clock(clock),
	.reset(reset)
);


// fifo_small_expand_key2_128_4_in_key
fifo_small #(
	.depth(64),
	.size(128)
) fifo_small_expand_key2_128_4_in_key(
	.datain(fifo_small_expand_key2_128_4_in_key_data),
	.dataout(expand_key2_128_4_in_key_data),
	.enr(expand_key2_128_4_in_key_rd),
	.enw(fifo_small_expand_key2_128_4_in_key_wr),
	.empty(expand_key2_128_4_in_key_empty),
	.full(fifo_small_expand_key2_128_4_in_key_full),
	
	// System Signal(s)
	.clk(clock),
	.rst(reset)
);

// actor expand_key2_128_4
expand_key2_128 actor_expand_key2_128_4 (
	// Input Signal(s)
	.in_key(expand_key2_128_4_in_key_data),
	.in_key_rd(expand_key2_128_4_in_key_rd),
	.in_key_empty(expand_key2_128_4_in_key_empty)
	,
	
	// Output Signal(s)
	.out_key(expand_key2_128_4_out_key_data),
	.out_key_wr(expand_key2_128_4_out_key_wr),
	.out_key_full(expand_key2_128_4_out_key_full)
		,
	
	// System Signal(s)
	.clock(clock),
	.reset(reset)
);


// fifo_small_expand_key3_128_4_in_key
fifo_small #(
	.depth(64),
	.size(128)
) fifo_small_expand_key3_128_4_in_key(
	.datain(fifo_small_expand_key3_128_4_in_key_data),
	.dataout(expand_key3_128_4_in_key_data),
	.enr(expand_key3_128_4_in_key_rd),
	.enw(fifo_small_expand_key3_128_4_in_key_wr),
	.empty(expand_key3_128_4_in_key_empty),
	.full(fifo_small_expand_key3_128_4_in_key_full),
	
	// System Signal(s)
	.clk(clock),
	.rst(reset)
);

// actor expand_key3_128_4
expand_key3_128 actor_expand_key3_128_4 (
	// Input Signal(s)
	.in_key(expand_key3_128_4_in_key_data),
	.in_key_rd(expand_key3_128_4_in_key_rd),
	.in_key_empty(expand_key3_128_4_in_key_empty)
	,
	
	// Output Signal(s)
	.out_key(expand_key3_128_4_out_key_data),
	.out_key_wr(expand_key3_128_4_out_key_wr),
	.out_key_full(expand_key3_128_4_out_key_full)
		,
	
	// System Signal(s)
	.clock(clock),
	.reset(reset)
);


// fifo_small_expand_key0_128_5_in_key
fifo_small #(
	.depth(64),
	.size(128)
) fifo_small_expand_key0_128_5_in_key(
	.datain(fifo_small_expand_key0_128_5_in_key_data),
	.dataout(expand_key0_128_5_in_key_data),
	.enr(expand_key0_128_5_in_key_rd),
	.enw(fifo_small_expand_key0_128_5_in_key_wr),
	.empty(expand_key0_128_5_in_key_empty),
	.full(fifo_small_expand_key0_128_5_in_key_full),
	
	// System Signal(s)
	.clk(clock),
	.rst(reset)
);
// fifo_small_expand_key0_128_5_in_rc
fifo_small #(
	.depth(64),
	.size(8)
) fifo_small_expand_key0_128_5_in_rc(
	.datain(fifo_small_expand_key0_128_5_in_rc_data),
	.dataout(expand_key0_128_5_in_rc_data),
	.enr(expand_key0_128_5_in_rc_rd),
	.enw(fifo_small_expand_key0_128_5_in_rc_wr),
	.empty(expand_key0_128_5_in_rc_empty),
	.full(fifo_small_expand_key0_128_5_in_rc_full),
	
	// System Signal(s)
	.clk(clock),
	.rst(reset)
);

// actor expand_key0_128_5
expand_key0_128 actor_expand_key0_128_5 (
	// Input Signal(s)
	.in_key(expand_key0_128_5_in_key_data),
	.in_key_rd(expand_key0_128_5_in_key_rd),
	.in_key_empty(expand_key0_128_5_in_key_empty),
	.in_rc(expand_key0_128_5_in_rc_data),
	.in_rc_rd(expand_key0_128_5_in_rc_rd),
	.in_rc_empty(expand_key0_128_5_in_rc_empty)
	,
	
	// Output Signal(s)
	.out_key(expand_key0_128_5_out_key_data),
	.out_key_wr(expand_key0_128_5_out_key_wr),
	.out_key_full(expand_key0_128_5_out_key_full)
		,
	
	// System Signal(s)
	.clock(clock),
	.reset(reset)
);


// fifo_small_expand_key1_128_5_in_key
fifo_small #(
	.depth(64),
	.size(128)
) fifo_small_expand_key1_128_5_in_key(
	.datain(fifo_small_expand_key1_128_5_in_key_data),
	.dataout(expand_key1_128_5_in_key_data),
	.enr(expand_key1_128_5_in_key_rd),
	.enw(fifo_small_expand_key1_128_5_in_key_wr),
	.empty(expand_key1_128_5_in_key_empty),
	.full(fifo_small_expand_key1_128_5_in_key_full),
	
	// System Signal(s)
	.clk(clock),
	.rst(reset)
);

// actor expand_key1_128_5
expand_key1_128 actor_expand_key1_128_5 (
	// Input Signal(s)
	.in_key(expand_key1_128_5_in_key_data),
	.in_key_rd(expand_key1_128_5_in_key_rd),
	.in_key_empty(expand_key1_128_5_in_key_empty)
	,
	
	// Output Signal(s)
	.out_key(expand_key1_128_5_out_key_data),
	.out_key_wr(expand_key1_128_5_out_key_wr),
	.out_key_full(expand_key1_128_5_out_key_full)
		,
	
	// System Signal(s)
	.clock(clock),
	.reset(reset)
);


// fifo_small_expand_key2_128_5_in_key
fifo_small #(
	.depth(64),
	.size(128)
) fifo_small_expand_key2_128_5_in_key(
	.datain(fifo_small_expand_key2_128_5_in_key_data),
	.dataout(expand_key2_128_5_in_key_data),
	.enr(expand_key2_128_5_in_key_rd),
	.enw(fifo_small_expand_key2_128_5_in_key_wr),
	.empty(expand_key2_128_5_in_key_empty),
	.full(fifo_small_expand_key2_128_5_in_key_full),
	
	// System Signal(s)
	.clk(clock),
	.rst(reset)
);

// actor expand_key2_128_5
expand_key2_128 actor_expand_key2_128_5 (
	// Input Signal(s)
	.in_key(expand_key2_128_5_in_key_data),
	.in_key_rd(expand_key2_128_5_in_key_rd),
	.in_key_empty(expand_key2_128_5_in_key_empty)
	,
	
	// Output Signal(s)
	.out_key(expand_key2_128_5_out_key_data),
	.out_key_wr(expand_key2_128_5_out_key_wr),
	.out_key_full(expand_key2_128_5_out_key_full)
		,
	
	// System Signal(s)
	.clock(clock),
	.reset(reset)
);


// fifo_small_expand_key3_128_5_in_key
fifo_small #(
	.depth(64),
	.size(128)
) fifo_small_expand_key3_128_5_in_key(
	.datain(fifo_small_expand_key3_128_5_in_key_data),
	.dataout(expand_key3_128_5_in_key_data),
	.enr(expand_key3_128_5_in_key_rd),
	.enw(fifo_small_expand_key3_128_5_in_key_wr),
	.empty(expand_key3_128_5_in_key_empty),
	.full(fifo_small_expand_key3_128_5_in_key_full),
	
	// System Signal(s)
	.clk(clock),
	.rst(reset)
);

// actor expand_key3_128_5
expand_key3_128 actor_expand_key3_128_5 (
	// Input Signal(s)
	.in_key(expand_key3_128_5_in_key_data),
	.in_key_rd(expand_key3_128_5_in_key_rd),
	.in_key_empty(expand_key3_128_5_in_key_empty)
	,
	
	// Output Signal(s)
	.out_key(expand_key3_128_5_out_key_data),
	.out_key_wr(expand_key3_128_5_out_key_wr),
	.out_key_full(expand_key3_128_5_out_key_full)
		,
	
	// System Signal(s)
	.clock(clock),
	.reset(reset)
);


// fifo_small_expand_key0_128_6_in_key
fifo_small #(
	.depth(64),
	.size(128)
) fifo_small_expand_key0_128_6_in_key(
	.datain(fifo_small_expand_key0_128_6_in_key_data),
	.dataout(expand_key0_128_6_in_key_data),
	.enr(expand_key0_128_6_in_key_rd),
	.enw(fifo_small_expand_key0_128_6_in_key_wr),
	.empty(expand_key0_128_6_in_key_empty),
	.full(fifo_small_expand_key0_128_6_in_key_full),
	
	// System Signal(s)
	.clk(clock),
	.rst(reset)
);
// fifo_small_expand_key0_128_6_in_rc
fifo_small #(
	.depth(64),
	.size(8)
) fifo_small_expand_key0_128_6_in_rc(
	.datain(fifo_small_expand_key0_128_6_in_rc_data),
	.dataout(expand_key0_128_6_in_rc_data),
	.enr(expand_key0_128_6_in_rc_rd),
	.enw(fifo_small_expand_key0_128_6_in_rc_wr),
	.empty(expand_key0_128_6_in_rc_empty),
	.full(fifo_small_expand_key0_128_6_in_rc_full),
	
	// System Signal(s)
	.clk(clock),
	.rst(reset)
);

// actor expand_key0_128_6
expand_key0_128 actor_expand_key0_128_6 (
	// Input Signal(s)
	.in_key(expand_key0_128_6_in_key_data),
	.in_key_rd(expand_key0_128_6_in_key_rd),
	.in_key_empty(expand_key0_128_6_in_key_empty),
	.in_rc(expand_key0_128_6_in_rc_data),
	.in_rc_rd(expand_key0_128_6_in_rc_rd),
	.in_rc_empty(expand_key0_128_6_in_rc_empty)
	,
	
	// Output Signal(s)
	.out_key(expand_key0_128_6_out_key_data),
	.out_key_wr(expand_key0_128_6_out_key_wr),
	.out_key_full(expand_key0_128_6_out_key_full)
		,
	
	// System Signal(s)
	.clock(clock),
	.reset(reset)
);


// fifo_small_expand_key1_128_6_in_key
fifo_small #(
	.depth(64),
	.size(128)
) fifo_small_expand_key1_128_6_in_key(
	.datain(fifo_small_expand_key1_128_6_in_key_data),
	.dataout(expand_key1_128_6_in_key_data),
	.enr(expand_key1_128_6_in_key_rd),
	.enw(fifo_small_expand_key1_128_6_in_key_wr),
	.empty(expand_key1_128_6_in_key_empty),
	.full(fifo_small_expand_key1_128_6_in_key_full),
	
	// System Signal(s)
	.clk(clock),
	.rst(reset)
);

// actor expand_key1_128_6
expand_key1_128 actor_expand_key1_128_6 (
	// Input Signal(s)
	.in_key(expand_key1_128_6_in_key_data),
	.in_key_rd(expand_key1_128_6_in_key_rd),
	.in_key_empty(expand_key1_128_6_in_key_empty)
	,
	
	// Output Signal(s)
	.out_key(expand_key1_128_6_out_key_data),
	.out_key_wr(expand_key1_128_6_out_key_wr),
	.out_key_full(expand_key1_128_6_out_key_full)
		,
	
	// System Signal(s)
	.clock(clock),
	.reset(reset)
);


// fifo_small_expand_key2_128_6_in_key
fifo_small #(
	.depth(64),
	.size(128)
) fifo_small_expand_key2_128_6_in_key(
	.datain(fifo_small_expand_key2_128_6_in_key_data),
	.dataout(expand_key2_128_6_in_key_data),
	.enr(expand_key2_128_6_in_key_rd),
	.enw(fifo_small_expand_key2_128_6_in_key_wr),
	.empty(expand_key2_128_6_in_key_empty),
	.full(fifo_small_expand_key2_128_6_in_key_full),
	
	// System Signal(s)
	.clk(clock),
	.rst(reset)
);

// actor expand_key2_128_6
expand_key2_128 actor_expand_key2_128_6 (
	// Input Signal(s)
	.in_key(expand_key2_128_6_in_key_data),
	.in_key_rd(expand_key2_128_6_in_key_rd),
	.in_key_empty(expand_key2_128_6_in_key_empty)
	,
	
	// Output Signal(s)
	.out_key(expand_key2_128_6_out_key_data),
	.out_key_wr(expand_key2_128_6_out_key_wr),
	.out_key_full(expand_key2_128_6_out_key_full)
		,
	
	// System Signal(s)
	.clock(clock),
	.reset(reset)
);


// fifo_small_expand_key3_128_6_in_key
fifo_small #(
	.depth(64),
	.size(128)
) fifo_small_expand_key3_128_6_in_key(
	.datain(fifo_small_expand_key3_128_6_in_key_data),
	.dataout(expand_key3_128_6_in_key_data),
	.enr(expand_key3_128_6_in_key_rd),
	.enw(fifo_small_expand_key3_128_6_in_key_wr),
	.empty(expand_key3_128_6_in_key_empty),
	.full(fifo_small_expand_key3_128_6_in_key_full),
	
	// System Signal(s)
	.clk(clock),
	.rst(reset)
);

// actor expand_key3_128_6
expand_key3_128 actor_expand_key3_128_6 (
	// Input Signal(s)
	.in_key(expand_key3_128_6_in_key_data),
	.in_key_rd(expand_key3_128_6_in_key_rd),
	.in_key_empty(expand_key3_128_6_in_key_empty)
	,
	
	// Output Signal(s)
	.out_key(expand_key3_128_6_out_key_data),
	.out_key_wr(expand_key3_128_6_out_key_wr),
	.out_key_full(expand_key3_128_6_out_key_full)
		,
	
	// System Signal(s)
	.clock(clock),
	.reset(reset)
);


// fifo_small_expand_key0_128_7_in_key
fifo_small #(
	.depth(64),
	.size(128)
) fifo_small_expand_key0_128_7_in_key(
	.datain(fifo_small_expand_key0_128_7_in_key_data),
	.dataout(expand_key0_128_7_in_key_data),
	.enr(expand_key0_128_7_in_key_rd),
	.enw(fifo_small_expand_key0_128_7_in_key_wr),
	.empty(expand_key0_128_7_in_key_empty),
	.full(fifo_small_expand_key0_128_7_in_key_full),
	
	// System Signal(s)
	.clk(clock),
	.rst(reset)
);
// fifo_small_expand_key0_128_7_in_rc
fifo_small #(
	.depth(64),
	.size(8)
) fifo_small_expand_key0_128_7_in_rc(
	.datain(fifo_small_expand_key0_128_7_in_rc_data),
	.dataout(expand_key0_128_7_in_rc_data),
	.enr(expand_key0_128_7_in_rc_rd),
	.enw(fifo_small_expand_key0_128_7_in_rc_wr),
	.empty(expand_key0_128_7_in_rc_empty),
	.full(fifo_small_expand_key0_128_7_in_rc_full),
	
	// System Signal(s)
	.clk(clock),
	.rst(reset)
);

// actor expand_key0_128_7
expand_key0_128 actor_expand_key0_128_7 (
	// Input Signal(s)
	.in_key(expand_key0_128_7_in_key_data),
	.in_key_rd(expand_key0_128_7_in_key_rd),
	.in_key_empty(expand_key0_128_7_in_key_empty),
	.in_rc(expand_key0_128_7_in_rc_data),
	.in_rc_rd(expand_key0_128_7_in_rc_rd),
	.in_rc_empty(expand_key0_128_7_in_rc_empty)
	,
	
	// Output Signal(s)
	.out_key(expand_key0_128_7_out_key_data),
	.out_key_wr(expand_key0_128_7_out_key_wr),
	.out_key_full(expand_key0_128_7_out_key_full)
		,
	
	// System Signal(s)
	.clock(clock),
	.reset(reset)
);


// fifo_small_expand_key1_128_7_in_key
fifo_small #(
	.depth(64),
	.size(128)
) fifo_small_expand_key1_128_7_in_key(
	.datain(fifo_small_expand_key1_128_7_in_key_data),
	.dataout(expand_key1_128_7_in_key_data),
	.enr(expand_key1_128_7_in_key_rd),
	.enw(fifo_small_expand_key1_128_7_in_key_wr),
	.empty(expand_key1_128_7_in_key_empty),
	.full(fifo_small_expand_key1_128_7_in_key_full),
	
	// System Signal(s)
	.clk(clock),
	.rst(reset)
);

// actor expand_key1_128_7
expand_key1_128 actor_expand_key1_128_7 (
	// Input Signal(s)
	.in_key(expand_key1_128_7_in_key_data),
	.in_key_rd(expand_key1_128_7_in_key_rd),
	.in_key_empty(expand_key1_128_7_in_key_empty)
	,
	
	// Output Signal(s)
	.out_key(expand_key1_128_7_out_key_data),
	.out_key_wr(expand_key1_128_7_out_key_wr),
	.out_key_full(expand_key1_128_7_out_key_full)
		,
	
	// System Signal(s)
	.clock(clock),
	.reset(reset)
);


// fifo_small_expand_key2_128_7_in_key
fifo_small #(
	.depth(64),
	.size(128)
) fifo_small_expand_key2_128_7_in_key(
	.datain(fifo_small_expand_key2_128_7_in_key_data),
	.dataout(expand_key2_128_7_in_key_data),
	.enr(expand_key2_128_7_in_key_rd),
	.enw(fifo_small_expand_key2_128_7_in_key_wr),
	.empty(expand_key2_128_7_in_key_empty),
	.full(fifo_small_expand_key2_128_7_in_key_full),
	
	// System Signal(s)
	.clk(clock),
	.rst(reset)
);

// actor expand_key2_128_7
expand_key2_128 actor_expand_key2_128_7 (
	// Input Signal(s)
	.in_key(expand_key2_128_7_in_key_data),
	.in_key_rd(expand_key2_128_7_in_key_rd),
	.in_key_empty(expand_key2_128_7_in_key_empty)
	,
	
	// Output Signal(s)
	.out_key(expand_key2_128_7_out_key_data),
	.out_key_wr(expand_key2_128_7_out_key_wr),
	.out_key_full(expand_key2_128_7_out_key_full)
		,
	
	// System Signal(s)
	.clock(clock),
	.reset(reset)
);


// fifo_small_expand_key3_128_7_in_key
fifo_small #(
	.depth(64),
	.size(128)
) fifo_small_expand_key3_128_7_in_key(
	.datain(fifo_small_expand_key3_128_7_in_key_data),
	.dataout(expand_key3_128_7_in_key_data),
	.enr(expand_key3_128_7_in_key_rd),
	.enw(fifo_small_expand_key3_128_7_in_key_wr),
	.empty(expand_key3_128_7_in_key_empty),
	.full(fifo_small_expand_key3_128_7_in_key_full),
	
	// System Signal(s)
	.clk(clock),
	.rst(reset)
);

// actor expand_key3_128_7
expand_key3_128 actor_expand_key3_128_7 (
	// Input Signal(s)
	.in_key(expand_key3_128_7_in_key_data),
	.in_key_rd(expand_key3_128_7_in_key_rd),
	.in_key_empty(expand_key3_128_7_in_key_empty)
	,
	
	// Output Signal(s)
	.out_key(expand_key3_128_7_out_key_data),
	.out_key_wr(expand_key3_128_7_out_key_wr),
	.out_key_full(expand_key3_128_7_out_key_full)
		,
	
	// System Signal(s)
	.clock(clock),
	.reset(reset)
);


// fifo_small_expand_key0_128_8_in_key
fifo_small #(
	.depth(64),
	.size(128)
) fifo_small_expand_key0_128_8_in_key(
	.datain(fifo_small_expand_key0_128_8_in_key_data),
	.dataout(expand_key0_128_8_in_key_data),
	.enr(expand_key0_128_8_in_key_rd),
	.enw(fifo_small_expand_key0_128_8_in_key_wr),
	.empty(expand_key0_128_8_in_key_empty),
	.full(fifo_small_expand_key0_128_8_in_key_full),
	
	// System Signal(s)
	.clk(clock),
	.rst(reset)
);
// fifo_small_expand_key0_128_8_in_rc
fifo_small #(
	.depth(64),
	.size(8)
) fifo_small_expand_key0_128_8_in_rc(
	.datain(fifo_small_expand_key0_128_8_in_rc_data),
	.dataout(expand_key0_128_8_in_rc_data),
	.enr(expand_key0_128_8_in_rc_rd),
	.enw(fifo_small_expand_key0_128_8_in_rc_wr),
	.empty(expand_key0_128_8_in_rc_empty),
	.full(fifo_small_expand_key0_128_8_in_rc_full),
	
	// System Signal(s)
	.clk(clock),
	.rst(reset)
);

// actor expand_key0_128_8
expand_key0_128 actor_expand_key0_128_8 (
	// Input Signal(s)
	.in_key(expand_key0_128_8_in_key_data),
	.in_key_rd(expand_key0_128_8_in_key_rd),
	.in_key_empty(expand_key0_128_8_in_key_empty),
	.in_rc(expand_key0_128_8_in_rc_data),
	.in_rc_rd(expand_key0_128_8_in_rc_rd),
	.in_rc_empty(expand_key0_128_8_in_rc_empty)
	,
	
	// Output Signal(s)
	.out_key(expand_key0_128_8_out_key_data),
	.out_key_wr(expand_key0_128_8_out_key_wr),
	.out_key_full(expand_key0_128_8_out_key_full)
		,
	
	// System Signal(s)
	.clock(clock),
	.reset(reset)
);


// fifo_small_expand_key1_128_8_in_key
fifo_small #(
	.depth(64),
	.size(128)
) fifo_small_expand_key1_128_8_in_key(
	.datain(fifo_small_expand_key1_128_8_in_key_data),
	.dataout(expand_key1_128_8_in_key_data),
	.enr(expand_key1_128_8_in_key_rd),
	.enw(fifo_small_expand_key1_128_8_in_key_wr),
	.empty(expand_key1_128_8_in_key_empty),
	.full(fifo_small_expand_key1_128_8_in_key_full),
	
	// System Signal(s)
	.clk(clock),
	.rst(reset)
);

// actor expand_key1_128_8
expand_key1_128 actor_expand_key1_128_8 (
	// Input Signal(s)
	.in_key(expand_key1_128_8_in_key_data),
	.in_key_rd(expand_key1_128_8_in_key_rd),
	.in_key_empty(expand_key1_128_8_in_key_empty)
	,
	
	// Output Signal(s)
	.out_key(expand_key1_128_8_out_key_data),
	.out_key_wr(expand_key1_128_8_out_key_wr),
	.out_key_full(expand_key1_128_8_out_key_full)
		,
	
	// System Signal(s)
	.clock(clock),
	.reset(reset)
);


// fifo_small_expand_key2_128_8_in_key
fifo_small #(
	.depth(64),
	.size(128)
) fifo_small_expand_key2_128_8_in_key(
	.datain(fifo_small_expand_key2_128_8_in_key_data),
	.dataout(expand_key2_128_8_in_key_data),
	.enr(expand_key2_128_8_in_key_rd),
	.enw(fifo_small_expand_key2_128_8_in_key_wr),
	.empty(expand_key2_128_8_in_key_empty),
	.full(fifo_small_expand_key2_128_8_in_key_full),
	
	// System Signal(s)
	.clk(clock),
	.rst(reset)
);

// actor expand_key2_128_8
expand_key2_128 actor_expand_key2_128_8 (
	// Input Signal(s)
	.in_key(expand_key2_128_8_in_key_data),
	.in_key_rd(expand_key2_128_8_in_key_rd),
	.in_key_empty(expand_key2_128_8_in_key_empty)
	,
	
	// Output Signal(s)
	.out_key(expand_key2_128_8_out_key_data),
	.out_key_wr(expand_key2_128_8_out_key_wr),
	.out_key_full(expand_key2_128_8_out_key_full)
		,
	
	// System Signal(s)
	.clock(clock),
	.reset(reset)
);


// fifo_small_expand_key3_128_8_in_key
fifo_small #(
	.depth(64),
	.size(128)
) fifo_small_expand_key3_128_8_in_key(
	.datain(fifo_small_expand_key3_128_8_in_key_data),
	.dataout(expand_key3_128_8_in_key_data),
	.enr(expand_key3_128_8_in_key_rd),
	.enw(fifo_small_expand_key3_128_8_in_key_wr),
	.empty(expand_key3_128_8_in_key_empty),
	.full(fifo_small_expand_key3_128_8_in_key_full),
	
	// System Signal(s)
	.clk(clock),
	.rst(reset)
);

// actor expand_key3_128_8
expand_key3_128 actor_expand_key3_128_8 (
	// Input Signal(s)
	.in_key(expand_key3_128_8_in_key_data),
	.in_key_rd(expand_key3_128_8_in_key_rd),
	.in_key_empty(expand_key3_128_8_in_key_empty)
	,
	
	// Output Signal(s)
	.out_key(expand_key3_128_8_out_key_data),
	.out_key_wr(expand_key3_128_8_out_key_wr),
	.out_key_full(expand_key3_128_8_out_key_full)
		,
	
	// System Signal(s)
	.clock(clock),
	.reset(reset)
);


// fifo_small_sub_bytes_9_in_state
fifo_small #(
	.depth(64),
	.size(128)
) fifo_small_sub_bytes_9_in_state(
	.datain(fifo_small_sub_bytes_9_in_state_data),
	.dataout(sub_bytes_9_in_state_data),
	.enr(sub_bytes_9_in_state_rd),
	.enw(fifo_small_sub_bytes_9_in_state_wr),
	.empty(sub_bytes_9_in_state_empty),
	.full(fifo_small_sub_bytes_9_in_state_full),
	
	// System Signal(s)
	.clk(clock),
	.rst(reset)
);

// actor sub_bytes_9
sub_bytes actor_sub_bytes_9 (
	// Input Signal(s)
	.in_state(sub_bytes_9_in_state_data),
	.in_state_rd(sub_bytes_9_in_state_rd),
	.in_state_empty(sub_bytes_9_in_state_empty)
	,
	
	// Output Signal(s)
	.out_state(sub_bytes_9_out_state_data),
	.out_state_wr(sub_bytes_9_out_state_wr),
	.out_state_full(sub_bytes_9_out_state_full)
		,
	
	// System Signal(s)
	.clock(clock),
	.reset(reset)
);


// fifo_small_shift_rows_9_in_state
fifo_small #(
	.depth(64),
	.size(128)
) fifo_small_shift_rows_9_in_state(
	.datain(fifo_small_shift_rows_9_in_state_data),
	.dataout(shift_rows_9_in_state_data),
	.enr(shift_rows_9_in_state_rd),
	.enw(fifo_small_shift_rows_9_in_state_wr),
	.empty(shift_rows_9_in_state_empty),
	.full(fifo_small_shift_rows_9_in_state_full),
	
	// System Signal(s)
	.clk(clock),
	.rst(reset)
);

// actor shift_rows_9
shift_rows actor_shift_rows_9 (
	// Input Signal(s)
	.in_state(shift_rows_9_in_state_data),
	.in_state_rd(shift_rows_9_in_state_rd),
	.in_state_empty(shift_rows_9_in_state_empty)
	,
	
	// Output Signal(s)
	.out_state(shift_rows_9_out_state_data),
	.out_state_wr(shift_rows_9_out_state_wr),
	.out_state_full(shift_rows_9_out_state_full)
		,
	
	// System Signal(s)
	.clock(clock),
	.reset(reset)
);


// fifo_small_mix_cols_8_in_state
fifo_small #(
	.depth(64),
	.size(128)
) fifo_small_mix_cols_8_in_state(
	.datain(fifo_small_mix_cols_8_in_state_data),
	.dataout(mix_cols_8_in_state_data),
	.enr(mix_cols_8_in_state_rd),
	.enw(fifo_small_mix_cols_8_in_state_wr),
	.empty(mix_cols_8_in_state_empty),
	.full(fifo_small_mix_cols_8_in_state_full),
	
	// System Signal(s)
	.clk(clock),
	.rst(reset)
);

// actor mix_cols_8
mix_cols actor_mix_cols_8 (
	// Input Signal(s)
	.in_state(mix_cols_8_in_state_data),
	.in_state_rd(mix_cols_8_in_state_rd),
	.in_state_empty(mix_cols_8_in_state_empty)
	,
	
	// Output Signal(s)
	.out_state(mix_cols_8_out_state_data),
	.out_state_wr(mix_cols_8_out_state_wr),
	.out_state_full(mix_cols_8_out_state_full)
		,
	
	// System Signal(s)
	.clock(clock),
	.reset(reset)
);


// fifo_small_add_round_key_10_in_state
fifo_small #(
	.depth(64),
	.size(128)
) fifo_small_add_round_key_10_in_state(
	.datain(fifo_small_add_round_key_10_in_state_data),
	.dataout(add_round_key_10_in_state_data),
	.enr(add_round_key_10_in_state_rd),
	.enw(fifo_small_add_round_key_10_in_state_wr),
	.empty(add_round_key_10_in_state_empty),
	.full(fifo_small_add_round_key_10_in_state_full),
	
	// System Signal(s)
	.clk(clock),
	.rst(reset)
);
// fifo_small_add_round_key_10_round_key
fifo_small #(
	.depth(64),
	.size(128)
) fifo_small_add_round_key_10_round_key(
	.datain(fifo_small_add_round_key_10_round_key_data),
	.dataout(add_round_key_10_round_key_data),
	.enr(add_round_key_10_round_key_rd),
	.enw(fifo_small_add_round_key_10_round_key_wr),
	.empty(add_round_key_10_round_key_empty),
	.full(fifo_small_add_round_key_10_round_key_full),
	
	// System Signal(s)
	.clk(clock),
	.rst(reset)
);

// actor add_round_key_10
add_round_key actor_add_round_key_10 (
	// Input Signal(s)
	.in_state(add_round_key_10_in_state_data),
	.in_state_rd(add_round_key_10_in_state_rd),
	.in_state_empty(add_round_key_10_in_state_empty),
	.round_key(add_round_key_10_round_key_data),
	.round_key_rd(add_round_key_10_round_key_rd),
	.round_key_empty(add_round_key_10_round_key_empty)
	,
	
	// Output Signal(s)
	.out_state(add_round_key_10_out_state_data),
	.out_state_wr(add_round_key_10_out_state_wr),
	.out_state_full(add_round_key_10_out_state_full)
		,
	
	// System Signal(s)
	.clock(clock),
	.reset(reset)
);


// fifo_small_expand_key0_128_9_in_key
fifo_small #(
	.depth(64),
	.size(128)
) fifo_small_expand_key0_128_9_in_key(
	.datain(fifo_small_expand_key0_128_9_in_key_data),
	.dataout(expand_key0_128_9_in_key_data),
	.enr(expand_key0_128_9_in_key_rd),
	.enw(fifo_small_expand_key0_128_9_in_key_wr),
	.empty(expand_key0_128_9_in_key_empty),
	.full(fifo_small_expand_key0_128_9_in_key_full),
	
	// System Signal(s)
	.clk(clock),
	.rst(reset)
);
// fifo_small_expand_key0_128_9_in_rc
fifo_small #(
	.depth(64),
	.size(8)
) fifo_small_expand_key0_128_9_in_rc(
	.datain(fifo_small_expand_key0_128_9_in_rc_data),
	.dataout(expand_key0_128_9_in_rc_data),
	.enr(expand_key0_128_9_in_rc_rd),
	.enw(fifo_small_expand_key0_128_9_in_rc_wr),
	.empty(expand_key0_128_9_in_rc_empty),
	.full(fifo_small_expand_key0_128_9_in_rc_full),
	
	// System Signal(s)
	.clk(clock),
	.rst(reset)
);

// actor expand_key0_128_9
expand_key0_128 actor_expand_key0_128_9 (
	// Input Signal(s)
	.in_key(expand_key0_128_9_in_key_data),
	.in_key_rd(expand_key0_128_9_in_key_rd),
	.in_key_empty(expand_key0_128_9_in_key_empty),
	.in_rc(expand_key0_128_9_in_rc_data),
	.in_rc_rd(expand_key0_128_9_in_rc_rd),
	.in_rc_empty(expand_key0_128_9_in_rc_empty)
	,
	
	// Output Signal(s)
	.out_key(expand_key0_128_9_out_key_data),
	.out_key_wr(expand_key0_128_9_out_key_wr),
	.out_key_full(expand_key0_128_9_out_key_full)
		,
	
	// System Signal(s)
	.clock(clock),
	.reset(reset)
);


// fifo_small_expand_key1_128_9_in_key
fifo_small #(
	.depth(64),
	.size(128)
) fifo_small_expand_key1_128_9_in_key(
	.datain(fifo_small_expand_key1_128_9_in_key_data),
	.dataout(expand_key1_128_9_in_key_data),
	.enr(expand_key1_128_9_in_key_rd),
	.enw(fifo_small_expand_key1_128_9_in_key_wr),
	.empty(expand_key1_128_9_in_key_empty),
	.full(fifo_small_expand_key1_128_9_in_key_full),
	
	// System Signal(s)
	.clk(clock),
	.rst(reset)
);

// actor expand_key1_128_9
expand_key1_128 actor_expand_key1_128_9 (
	// Input Signal(s)
	.in_key(expand_key1_128_9_in_key_data),
	.in_key_rd(expand_key1_128_9_in_key_rd),
	.in_key_empty(expand_key1_128_9_in_key_empty)
	,
	
	// Output Signal(s)
	.out_key(expand_key1_128_9_out_key_data),
	.out_key_wr(expand_key1_128_9_out_key_wr),
	.out_key_full(expand_key1_128_9_out_key_full)
		,
	
	// System Signal(s)
	.clock(clock),
	.reset(reset)
);


// fifo_small_expand_key2_128_9_in_key
fifo_small #(
	.depth(64),
	.size(128)
) fifo_small_expand_key2_128_9_in_key(
	.datain(fifo_small_expand_key2_128_9_in_key_data),
	.dataout(expand_key2_128_9_in_key_data),
	.enr(expand_key2_128_9_in_key_rd),
	.enw(fifo_small_expand_key2_128_9_in_key_wr),
	.empty(expand_key2_128_9_in_key_empty),
	.full(fifo_small_expand_key2_128_9_in_key_full),
	
	// System Signal(s)
	.clk(clock),
	.rst(reset)
);

// actor expand_key2_128_9
expand_key2_128 actor_expand_key2_128_9 (
	// Input Signal(s)
	.in_key(expand_key2_128_9_in_key_data),
	.in_key_rd(expand_key2_128_9_in_key_rd),
	.in_key_empty(expand_key2_128_9_in_key_empty)
	,
	
	// Output Signal(s)
	.out_key(expand_key2_128_9_out_key_data),
	.out_key_wr(expand_key2_128_9_out_key_wr),
	.out_key_full(expand_key2_128_9_out_key_full)
		,
	
	// System Signal(s)
	.clock(clock),
	.reset(reset)
);


// fifo_small_expand_key3_128_9_in_key
fifo_small #(
	.depth(64),
	.size(128)
) fifo_small_expand_key3_128_9_in_key(
	.datain(fifo_small_expand_key3_128_9_in_key_data),
	.dataout(expand_key3_128_9_in_key_data),
	.enr(expand_key3_128_9_in_key_rd),
	.enw(fifo_small_expand_key3_128_9_in_key_wr),
	.empty(expand_key3_128_9_in_key_empty),
	.full(fifo_small_expand_key3_128_9_in_key_full),
	
	// System Signal(s)
	.clk(clock),
	.rst(reset)
);

// actor expand_key3_128_9
expand_key3_128 actor_expand_key3_128_9 (
	// Input Signal(s)
	.in_key(expand_key3_128_9_in_key_data),
	.in_key_rd(expand_key3_128_9_in_key_rd),
	.in_key_empty(expand_key3_128_9_in_key_empty)
	,
	
	// Output Signal(s)
	.out_key(expand_key3_128_9_out_key_data),
	.out_key_wr(expand_key3_128_9_out_key_wr),
	.out_key_full(expand_key3_128_9_out_key_full)
		,
	
	// System Signal(s)
	.clock(clock),
	.reset(reset)
);


// Module(s) Assignments
assign fifo_small_read8x16_1_in_token_data = text_data;
assign fifo_small_read8x16_1_in_token_wr = text_wr;
assign text_full = fifo_small_read8x16_1_in_token_full;

assign fifo_small_read8x16_0_in_token_data = key_data;
assign fifo_small_read8x16_0_in_token_wr = key_wr;
assign key_full = fifo_small_read8x16_0_in_token_full;

assign fifo_small_expand_key0_128_0_in_key_data = read8x16_0_out_token_data;
assign fifo_small_expand_key0_128_0_in_key_wr = read8x16_0_out_token_wr;
assign read8x16_0_out_token_full =
fifo_small_expand_key0_128_0_in_key_full || 
fifo_small_add_round_key_0_round_key_full 
;

assign fifo_small_expand_key0_128_0_in_rc_data = rc_data;
assign fifo_small_expand_key0_128_0_in_rc_wr = rc_wr;
assign rc_full =		
fifo_small_expand_key0_128_0_in_rc_full || 
fifo_small_expand_key0_128_1_in_rc_full || 
fifo_small_expand_key0_128_2_in_rc_full || 
fifo_small_expand_key0_128_3_in_rc_full || 
fifo_small_expand_key0_128_4_in_rc_full || 
fifo_small_expand_key0_128_5_in_rc_full || 
fifo_small_expand_key0_128_6_in_rc_full || 
fifo_small_expand_key0_128_7_in_rc_full || 
fifo_small_expand_key0_128_8_in_rc_full || 
fifo_small_expand_key0_128_9_in_rc_full 
;

assign fifo_small_expand_key0_128_1_in_rc_data = rc_data;
assign fifo_small_expand_key0_128_1_in_rc_wr = rc_wr;

assign fifo_small_expand_key0_128_1_in_key_data = expand_key3_128_0_out_key_data;
assign fifo_small_expand_key0_128_1_in_key_wr = expand_key3_128_0_out_key_wr;
assign expand_key3_128_0_out_key_full =
fifo_small_expand_key0_128_1_in_key_full || 
fifo_small_add_round_key_2_round_key_full 
;

assign fifo_small_expand_key0_128_2_in_rc_data = rc_data;
assign fifo_small_expand_key0_128_2_in_rc_wr = rc_wr;

assign fifo_small_expand_key0_128_2_in_key_data = expand_key3_128_1_out_key_data;
assign fifo_small_expand_key0_128_2_in_key_wr = expand_key3_128_1_out_key_wr;
assign expand_key3_128_1_out_key_full =
fifo_small_expand_key0_128_2_in_key_full || 
fifo_small_add_round_key_3_round_key_full 
;

assign fifo_small_expand_key0_128_3_in_rc_data = rc_data;
assign fifo_small_expand_key0_128_3_in_rc_wr = rc_wr;

assign fifo_small_expand_key0_128_3_in_key_data = expand_key3_128_2_out_key_data;
assign fifo_small_expand_key0_128_3_in_key_wr = expand_key3_128_2_out_key_wr;
assign expand_key3_128_2_out_key_full =
fifo_small_expand_key0_128_3_in_key_full || 
fifo_small_add_round_key_4_round_key_full 
;

assign fifo_small_expand_key0_128_4_in_rc_data = rc_data;
assign fifo_small_expand_key0_128_4_in_rc_wr = rc_wr;

assign fifo_small_expand_key0_128_4_in_key_data = expand_key3_128_3_out_key_data;
assign fifo_small_expand_key0_128_4_in_key_wr = expand_key3_128_3_out_key_wr;
assign expand_key3_128_3_out_key_full =
fifo_small_expand_key0_128_4_in_key_full || 
fifo_small_add_round_key_5_round_key_full 
;

assign fifo_small_expand_key0_128_5_in_rc_data = rc_data;
assign fifo_small_expand_key0_128_5_in_rc_wr = rc_wr;

assign fifo_small_expand_key0_128_5_in_key_data = expand_key3_128_4_out_key_data;
assign fifo_small_expand_key0_128_5_in_key_wr = expand_key3_128_4_out_key_wr;
assign expand_key3_128_4_out_key_full =
fifo_small_expand_key0_128_5_in_key_full || 
fifo_small_add_round_key_6_round_key_full 
;

assign fifo_small_expand_key0_128_6_in_rc_data = rc_data;
assign fifo_small_expand_key0_128_6_in_rc_wr = rc_wr;

assign fifo_small_expand_key0_128_6_in_key_data = expand_key3_128_5_out_key_data;
assign fifo_small_expand_key0_128_6_in_key_wr = expand_key3_128_5_out_key_wr;
assign expand_key3_128_5_out_key_full =
fifo_small_expand_key0_128_6_in_key_full || 
fifo_small_add_round_key_7_round_key_full 
;

assign fifo_small_expand_key0_128_7_in_rc_data = rc_data;
assign fifo_small_expand_key0_128_7_in_rc_wr = rc_wr;

assign fifo_small_expand_key0_128_7_in_key_data = expand_key3_128_6_out_key_data;
assign fifo_small_expand_key0_128_7_in_key_wr = expand_key3_128_6_out_key_wr;
assign expand_key3_128_6_out_key_full =
fifo_small_expand_key0_128_7_in_key_full || 
fifo_small_add_round_key_8_round_key_full 
;

assign fifo_small_expand_key0_128_8_in_rc_data = rc_data;
assign fifo_small_expand_key0_128_8_in_rc_wr = rc_wr;

assign fifo_small_expand_key0_128_8_in_key_data = expand_key3_128_7_out_key_data;
assign fifo_small_expand_key0_128_8_in_key_wr = expand_key3_128_7_out_key_wr;
assign expand_key3_128_7_out_key_full =
fifo_small_expand_key0_128_8_in_key_full || 
fifo_small_add_round_key_9_round_key_full 
;

assign fifo_small_expand_key0_128_9_in_rc_data = rc_data;
assign fifo_small_expand_key0_128_9_in_rc_wr = rc_wr;

assign fifo_small_expand_key0_128_9_in_key_data = expand_key3_128_8_out_key_data;
assign fifo_small_expand_key0_128_9_in_key_wr = expand_key3_128_8_out_key_wr;
assign expand_key3_128_8_out_key_full =
fifo_small_expand_key0_128_9_in_key_full || 
fifo_small_add_round_key_10_round_key_full 
;

assign fifo_small_add_round_key_0_in_state_data = read8x16_1_out_token_data;
assign fifo_small_add_round_key_0_in_state_wr = read8x16_1_out_token_wr;
assign read8x16_1_out_token_full = fifo_small_add_round_key_0_in_state_full;

assign fifo_small_add_round_key_0_round_key_data = read8x16_0_out_token_data;
assign fifo_small_add_round_key_0_round_key_wr = read8x16_0_out_token_wr;

assign fifo_small_expand_key1_128_0_in_key_data = expand_key0_128_0_out_key_data;
assign fifo_small_expand_key1_128_0_in_key_wr = expand_key0_128_0_out_key_wr;
assign expand_key0_128_0_out_key_full = fifo_small_expand_key1_128_0_in_key_full;

assign fifo_small_expand_key1_128_1_in_key_data = expand_key0_128_1_out_key_data;
assign fifo_small_expand_key1_128_1_in_key_wr = expand_key0_128_1_out_key_wr;
assign expand_key0_128_1_out_key_full = fifo_small_expand_key1_128_1_in_key_full;

assign fifo_small_expand_key1_128_2_in_key_data = expand_key0_128_2_out_key_data;
assign fifo_small_expand_key1_128_2_in_key_wr = expand_key0_128_2_out_key_wr;
assign expand_key0_128_2_out_key_full = fifo_small_expand_key1_128_2_in_key_full;

assign fifo_small_expand_key1_128_3_in_key_data = expand_key0_128_3_out_key_data;
assign fifo_small_expand_key1_128_3_in_key_wr = expand_key0_128_3_out_key_wr;
assign expand_key0_128_3_out_key_full = fifo_small_expand_key1_128_3_in_key_full;

assign fifo_small_expand_key1_128_4_in_key_data = expand_key0_128_4_out_key_data;
assign fifo_small_expand_key1_128_4_in_key_wr = expand_key0_128_4_out_key_wr;
assign expand_key0_128_4_out_key_full = fifo_small_expand_key1_128_4_in_key_full;

assign fifo_small_expand_key1_128_5_in_key_data = expand_key0_128_5_out_key_data;
assign fifo_small_expand_key1_128_5_in_key_wr = expand_key0_128_5_out_key_wr;
assign expand_key0_128_5_out_key_full = fifo_small_expand_key1_128_5_in_key_full;

assign fifo_small_expand_key1_128_6_in_key_data = expand_key0_128_6_out_key_data;
assign fifo_small_expand_key1_128_6_in_key_wr = expand_key0_128_6_out_key_wr;
assign expand_key0_128_6_out_key_full = fifo_small_expand_key1_128_6_in_key_full;

assign fifo_small_expand_key1_128_7_in_key_data = expand_key0_128_7_out_key_data;
assign fifo_small_expand_key1_128_7_in_key_wr = expand_key0_128_7_out_key_wr;
assign expand_key0_128_7_out_key_full = fifo_small_expand_key1_128_7_in_key_full;

assign fifo_small_expand_key1_128_8_in_key_data = expand_key0_128_8_out_key_data;
assign fifo_small_expand_key1_128_8_in_key_wr = expand_key0_128_8_out_key_wr;
assign expand_key0_128_8_out_key_full = fifo_small_expand_key1_128_8_in_key_full;

assign fifo_small_expand_key1_128_9_in_key_data = expand_key0_128_9_out_key_data;
assign fifo_small_expand_key1_128_9_in_key_wr = expand_key0_128_9_out_key_wr;
assign expand_key0_128_9_out_key_full = fifo_small_expand_key1_128_9_in_key_full;

assign fifo_small_sub_bytes_1_in_state_data = add_round_key_0_out_state_data;
assign fifo_small_sub_bytes_1_in_state_wr = add_round_key_0_out_state_wr;
assign add_round_key_0_out_state_full = fifo_small_sub_bytes_1_in_state_full;

assign fifo_small_expand_key2_128_0_in_key_data = expand_key1_128_0_out_key_data;
assign fifo_small_expand_key2_128_0_in_key_wr = expand_key1_128_0_out_key_wr;
assign expand_key1_128_0_out_key_full = fifo_small_expand_key2_128_0_in_key_full;

assign fifo_small_expand_key2_128_1_in_key_data = expand_key1_128_1_out_key_data;
assign fifo_small_expand_key2_128_1_in_key_wr = expand_key1_128_1_out_key_wr;
assign expand_key1_128_1_out_key_full = fifo_small_expand_key2_128_1_in_key_full;

assign fifo_small_expand_key2_128_2_in_key_data = expand_key1_128_2_out_key_data;
assign fifo_small_expand_key2_128_2_in_key_wr = expand_key1_128_2_out_key_wr;
assign expand_key1_128_2_out_key_full = fifo_small_expand_key2_128_2_in_key_full;

assign fifo_small_expand_key2_128_3_in_key_data = expand_key1_128_3_out_key_data;
assign fifo_small_expand_key2_128_3_in_key_wr = expand_key1_128_3_out_key_wr;
assign expand_key1_128_3_out_key_full = fifo_small_expand_key2_128_3_in_key_full;

assign fifo_small_expand_key2_128_4_in_key_data = expand_key1_128_4_out_key_data;
assign fifo_small_expand_key2_128_4_in_key_wr = expand_key1_128_4_out_key_wr;
assign expand_key1_128_4_out_key_full = fifo_small_expand_key2_128_4_in_key_full;

assign fifo_small_expand_key2_128_5_in_key_data = expand_key1_128_5_out_key_data;
assign fifo_small_expand_key2_128_5_in_key_wr = expand_key1_128_5_out_key_wr;
assign expand_key1_128_5_out_key_full = fifo_small_expand_key2_128_5_in_key_full;

assign fifo_small_expand_key2_128_6_in_key_data = expand_key1_128_6_out_key_data;
assign fifo_small_expand_key2_128_6_in_key_wr = expand_key1_128_6_out_key_wr;
assign expand_key1_128_6_out_key_full = fifo_small_expand_key2_128_6_in_key_full;

assign fifo_small_expand_key2_128_7_in_key_data = expand_key1_128_7_out_key_data;
assign fifo_small_expand_key2_128_7_in_key_wr = expand_key1_128_7_out_key_wr;
assign expand_key1_128_7_out_key_full = fifo_small_expand_key2_128_7_in_key_full;

assign fifo_small_expand_key2_128_8_in_key_data = expand_key1_128_8_out_key_data;
assign fifo_small_expand_key2_128_8_in_key_wr = expand_key1_128_8_out_key_wr;
assign expand_key1_128_8_out_key_full = fifo_small_expand_key2_128_8_in_key_full;

assign fifo_small_expand_key2_128_9_in_key_data = expand_key1_128_9_out_key_data;
assign fifo_small_expand_key2_128_9_in_key_wr = expand_key1_128_9_out_key_wr;
assign expand_key1_128_9_out_key_full = fifo_small_expand_key2_128_9_in_key_full;

assign fifo_small_shift_rows_1_in_state_data = sub_bytes_1_out_state_data;
assign fifo_small_shift_rows_1_in_state_wr = sub_bytes_1_out_state_wr;
assign sub_bytes_1_out_state_full = fifo_small_shift_rows_1_in_state_full;

assign fifo_small_expand_key3_128_0_in_key_data = expand_key2_128_0_out_key_data;
assign fifo_small_expand_key3_128_0_in_key_wr = expand_key2_128_0_out_key_wr;
assign expand_key2_128_0_out_key_full = fifo_small_expand_key3_128_0_in_key_full;

assign fifo_small_expand_key3_128_1_in_key_data = expand_key2_128_1_out_key_data;
assign fifo_small_expand_key3_128_1_in_key_wr = expand_key2_128_1_out_key_wr;
assign expand_key2_128_1_out_key_full = fifo_small_expand_key3_128_1_in_key_full;

assign fifo_small_expand_key3_128_2_in_key_data = expand_key2_128_2_out_key_data;
assign fifo_small_expand_key3_128_2_in_key_wr = expand_key2_128_2_out_key_wr;
assign expand_key2_128_2_out_key_full = fifo_small_expand_key3_128_2_in_key_full;

assign fifo_small_expand_key3_128_3_in_key_data = expand_key2_128_3_out_key_data;
assign fifo_small_expand_key3_128_3_in_key_wr = expand_key2_128_3_out_key_wr;
assign expand_key2_128_3_out_key_full = fifo_small_expand_key3_128_3_in_key_full;

assign fifo_small_expand_key3_128_4_in_key_data = expand_key2_128_4_out_key_data;
assign fifo_small_expand_key3_128_4_in_key_wr = expand_key2_128_4_out_key_wr;
assign expand_key2_128_4_out_key_full = fifo_small_expand_key3_128_4_in_key_full;

assign fifo_small_expand_key3_128_5_in_key_data = expand_key2_128_5_out_key_data;
assign fifo_small_expand_key3_128_5_in_key_wr = expand_key2_128_5_out_key_wr;
assign expand_key2_128_5_out_key_full = fifo_small_expand_key3_128_5_in_key_full;

assign fifo_small_expand_key3_128_6_in_key_data = expand_key2_128_6_out_key_data;
assign fifo_small_expand_key3_128_6_in_key_wr = expand_key2_128_6_out_key_wr;
assign expand_key2_128_6_out_key_full = fifo_small_expand_key3_128_6_in_key_full;

assign fifo_small_expand_key3_128_7_in_key_data = expand_key2_128_7_out_key_data;
assign fifo_small_expand_key3_128_7_in_key_wr = expand_key2_128_7_out_key_wr;
assign expand_key2_128_7_out_key_full = fifo_small_expand_key3_128_7_in_key_full;

assign fifo_small_expand_key3_128_8_in_key_data = expand_key2_128_8_out_key_data;
assign fifo_small_expand_key3_128_8_in_key_wr = expand_key2_128_8_out_key_wr;
assign expand_key2_128_8_out_key_full = fifo_small_expand_key3_128_8_in_key_full;

assign fifo_small_expand_key3_128_9_in_key_data = expand_key2_128_9_out_key_data;
assign fifo_small_expand_key3_128_9_in_key_wr = expand_key2_128_9_out_key_wr;
assign expand_key2_128_9_out_key_full = fifo_small_expand_key3_128_9_in_key_full;

assign fifo_small_mix_cols_0_in_state_data = shift_rows_1_out_state_data;
assign fifo_small_mix_cols_0_in_state_wr = shift_rows_1_out_state_wr;
assign shift_rows_1_out_state_full = fifo_small_mix_cols_0_in_state_full;

assign fifo_small_add_round_key_2_in_state_data = mix_cols_0_out_state_data;
assign fifo_small_add_round_key_2_in_state_wr = mix_cols_0_out_state_wr;
assign mix_cols_0_out_state_full = fifo_small_add_round_key_2_in_state_full;

assign fifo_small_add_round_key_2_round_key_data = expand_key3_128_0_out_key_data;
assign fifo_small_add_round_key_2_round_key_wr = expand_key3_128_0_out_key_wr;

assign fifo_small_add_round_key_3_in_state_data = mix_cols_1_out_state_data;
assign fifo_small_add_round_key_3_in_state_wr = mix_cols_1_out_state_wr;
assign mix_cols_1_out_state_full = fifo_small_add_round_key_3_in_state_full;

assign fifo_small_add_round_key_3_round_key_data = expand_key3_128_1_out_key_data;
assign fifo_small_add_round_key_3_round_key_wr = expand_key3_128_1_out_key_wr;

assign fifo_small_add_round_key_4_in_state_data = mix_cols_2_out_state_data;
assign fifo_small_add_round_key_4_in_state_wr = mix_cols_2_out_state_wr;
assign mix_cols_2_out_state_full = fifo_small_add_round_key_4_in_state_full;

assign fifo_small_add_round_key_4_round_key_data = expand_key3_128_2_out_key_data;
assign fifo_small_add_round_key_4_round_key_wr = expand_key3_128_2_out_key_wr;

assign fifo_small_add_round_key_5_in_state_data = mix_cols_3_out_state_data;
assign fifo_small_add_round_key_5_in_state_wr = mix_cols_3_out_state_wr;
assign mix_cols_3_out_state_full = fifo_small_add_round_key_5_in_state_full;

assign fifo_small_add_round_key_5_round_key_data = expand_key3_128_3_out_key_data;
assign fifo_small_add_round_key_5_round_key_wr = expand_key3_128_3_out_key_wr;

assign fifo_small_add_round_key_6_in_state_data = mix_cols_4_out_state_data;
assign fifo_small_add_round_key_6_in_state_wr = mix_cols_4_out_state_wr;
assign mix_cols_4_out_state_full = fifo_small_add_round_key_6_in_state_full;

assign fifo_small_add_round_key_6_round_key_data = expand_key3_128_4_out_key_data;
assign fifo_small_add_round_key_6_round_key_wr = expand_key3_128_4_out_key_wr;

assign fifo_small_add_round_key_7_in_state_data = mix_cols_5_out_state_data;
assign fifo_small_add_round_key_7_in_state_wr = mix_cols_5_out_state_wr;
assign mix_cols_5_out_state_full = fifo_small_add_round_key_7_in_state_full;

assign fifo_small_add_round_key_7_round_key_data = expand_key3_128_5_out_key_data;
assign fifo_small_add_round_key_7_round_key_wr = expand_key3_128_5_out_key_wr;

assign fifo_small_add_round_key_8_in_state_data = mix_cols_6_out_state_data;
assign fifo_small_add_round_key_8_in_state_wr = mix_cols_6_out_state_wr;
assign mix_cols_6_out_state_full = fifo_small_add_round_key_8_in_state_full;

assign fifo_small_add_round_key_8_round_key_data = expand_key3_128_6_out_key_data;
assign fifo_small_add_round_key_8_round_key_wr = expand_key3_128_6_out_key_wr;

assign fifo_small_add_round_key_9_in_state_data = mix_cols_7_out_state_data;
assign fifo_small_add_round_key_9_in_state_wr = mix_cols_7_out_state_wr;
assign mix_cols_7_out_state_full = fifo_small_add_round_key_9_in_state_full;

assign fifo_small_add_round_key_9_round_key_data = expand_key3_128_7_out_key_data;
assign fifo_small_add_round_key_9_round_key_wr = expand_key3_128_7_out_key_wr;

assign fifo_small_add_round_key_10_in_state_data = mix_cols_8_out_state_data;
assign fifo_small_add_round_key_10_in_state_wr = mix_cols_8_out_state_wr;
assign mix_cols_8_out_state_full = fifo_small_add_round_key_10_in_state_full;

assign fifo_small_add_round_key_10_round_key_data = expand_key3_128_8_out_key_data;
assign fifo_small_add_round_key_10_round_key_wr = expand_key3_128_8_out_key_wr;

assign fifo_small_add_round_key_1_in_state_data = shift_rows_0_out_state_data;
assign fifo_small_add_round_key_1_in_state_wr = shift_rows_0_out_state_wr;
assign shift_rows_0_out_state_full = fifo_small_add_round_key_1_in_state_full;

assign fifo_small_add_round_key_1_round_key_data = expand_key3_128_9_out_key_data;
assign fifo_small_add_round_key_1_round_key_wr = expand_key3_128_9_out_key_wr;
assign expand_key3_128_9_out_key_full = fifo_small_add_round_key_1_round_key_full;

assign fifo_small_sub_bytes_2_in_state_data = add_round_key_2_out_state_data;
assign fifo_small_sub_bytes_2_in_state_wr = add_round_key_2_out_state_wr;
assign add_round_key_2_out_state_full = fifo_small_sub_bytes_2_in_state_full;

assign fifo_small_sub_bytes_3_in_state_data = add_round_key_3_out_state_data;
assign fifo_small_sub_bytes_3_in_state_wr = add_round_key_3_out_state_wr;
assign add_round_key_3_out_state_full = fifo_small_sub_bytes_3_in_state_full;

assign fifo_small_sub_bytes_4_in_state_data = add_round_key_4_out_state_data;
assign fifo_small_sub_bytes_4_in_state_wr = add_round_key_4_out_state_wr;
assign add_round_key_4_out_state_full = fifo_small_sub_bytes_4_in_state_full;

assign fifo_small_sub_bytes_5_in_state_data = add_round_key_5_out_state_data;
assign fifo_small_sub_bytes_5_in_state_wr = add_round_key_5_out_state_wr;
assign add_round_key_5_out_state_full = fifo_small_sub_bytes_5_in_state_full;

assign fifo_small_sub_bytes_6_in_state_data = add_round_key_6_out_state_data;
assign fifo_small_sub_bytes_6_in_state_wr = add_round_key_6_out_state_wr;
assign add_round_key_6_out_state_full = fifo_small_sub_bytes_6_in_state_full;

assign fifo_small_sub_bytes_7_in_state_data = add_round_key_7_out_state_data;
assign fifo_small_sub_bytes_7_in_state_wr = add_round_key_7_out_state_wr;
assign add_round_key_7_out_state_full = fifo_small_sub_bytes_7_in_state_full;

assign fifo_small_sub_bytes_8_in_state_data = add_round_key_8_out_state_data;
assign fifo_small_sub_bytes_8_in_state_wr = add_round_key_8_out_state_wr;
assign add_round_key_8_out_state_full = fifo_small_sub_bytes_8_in_state_full;

assign fifo_small_sub_bytes_9_in_state_data = add_round_key_9_out_state_data;
assign fifo_small_sub_bytes_9_in_state_wr = add_round_key_9_out_state_wr;
assign add_round_key_9_out_state_full = fifo_small_sub_bytes_9_in_state_full;

assign fifo_small_sub_bytes_0_in_state_data = add_round_key_10_out_state_data;
assign fifo_small_sub_bytes_0_in_state_wr = add_round_key_10_out_state_wr;
assign add_round_key_10_out_state_full = fifo_small_sub_bytes_0_in_state_full;

assign fifo_small_write16x8_0_in_token_data = add_round_key_1_out_state_data;
assign fifo_small_write16x8_0_in_token_wr = add_round_key_1_out_state_wr;
assign add_round_key_1_out_state_full = fifo_small_write16x8_0_in_token_full;

assign fifo_small_shift_rows_2_in_state_data = sub_bytes_2_out_state_data;
assign fifo_small_shift_rows_2_in_state_wr = sub_bytes_2_out_state_wr;
assign sub_bytes_2_out_state_full = fifo_small_shift_rows_2_in_state_full;

assign fifo_small_shift_rows_3_in_state_data = sub_bytes_3_out_state_data;
assign fifo_small_shift_rows_3_in_state_wr = sub_bytes_3_out_state_wr;
assign sub_bytes_3_out_state_full = fifo_small_shift_rows_3_in_state_full;

assign fifo_small_shift_rows_4_in_state_data = sub_bytes_4_out_state_data;
assign fifo_small_shift_rows_4_in_state_wr = sub_bytes_4_out_state_wr;
assign sub_bytes_4_out_state_full = fifo_small_shift_rows_4_in_state_full;

assign fifo_small_shift_rows_5_in_state_data = sub_bytes_5_out_state_data;
assign fifo_small_shift_rows_5_in_state_wr = sub_bytes_5_out_state_wr;
assign sub_bytes_5_out_state_full = fifo_small_shift_rows_5_in_state_full;

assign fifo_small_shift_rows_6_in_state_data = sub_bytes_6_out_state_data;
assign fifo_small_shift_rows_6_in_state_wr = sub_bytes_6_out_state_wr;
assign sub_bytes_6_out_state_full = fifo_small_shift_rows_6_in_state_full;

assign fifo_small_shift_rows_7_in_state_data = sub_bytes_7_out_state_data;
assign fifo_small_shift_rows_7_in_state_wr = sub_bytes_7_out_state_wr;
assign sub_bytes_7_out_state_full = fifo_small_shift_rows_7_in_state_full;

assign fifo_small_shift_rows_8_in_state_data = sub_bytes_8_out_state_data;
assign fifo_small_shift_rows_8_in_state_wr = sub_bytes_8_out_state_wr;
assign sub_bytes_8_out_state_full = fifo_small_shift_rows_8_in_state_full;

assign fifo_small_shift_rows_9_in_state_data = sub_bytes_9_out_state_data;
assign fifo_small_shift_rows_9_in_state_wr = sub_bytes_9_out_state_wr;
assign sub_bytes_9_out_state_full = fifo_small_shift_rows_9_in_state_full;

assign fifo_small_shift_rows_0_in_state_data = sub_bytes_0_out_state_data;
assign fifo_small_shift_rows_0_in_state_wr = sub_bytes_0_out_state_wr;
assign sub_bytes_0_out_state_full = fifo_small_shift_rows_0_in_state_full;

assign chiped_text_data = write16x8_0_out_token_data;
assign chiped_text_wr = write16x8_0_out_token_wr;
assign write16x8_0_out_token_full = chiped_text_full;

assign fifo_small_mix_cols_1_in_state_data = shift_rows_2_out_state_data;
assign fifo_small_mix_cols_1_in_state_wr = shift_rows_2_out_state_wr;
assign shift_rows_2_out_state_full = fifo_small_mix_cols_1_in_state_full;

assign fifo_small_mix_cols_2_in_state_data = shift_rows_3_out_state_data;
assign fifo_small_mix_cols_2_in_state_wr = shift_rows_3_out_state_wr;
assign shift_rows_3_out_state_full = fifo_small_mix_cols_2_in_state_full;

assign fifo_small_mix_cols_3_in_state_data = shift_rows_4_out_state_data;
assign fifo_small_mix_cols_3_in_state_wr = shift_rows_4_out_state_wr;
assign shift_rows_4_out_state_full = fifo_small_mix_cols_3_in_state_full;

assign fifo_small_mix_cols_4_in_state_data = shift_rows_5_out_state_data;
assign fifo_small_mix_cols_4_in_state_wr = shift_rows_5_out_state_wr;
assign shift_rows_5_out_state_full = fifo_small_mix_cols_4_in_state_full;

assign fifo_small_mix_cols_5_in_state_data = shift_rows_6_out_state_data;
assign fifo_small_mix_cols_5_in_state_wr = shift_rows_6_out_state_wr;
assign shift_rows_6_out_state_full = fifo_small_mix_cols_5_in_state_full;

assign fifo_small_mix_cols_6_in_state_data = shift_rows_7_out_state_data;
assign fifo_small_mix_cols_6_in_state_wr = shift_rows_7_out_state_wr;
assign shift_rows_7_out_state_full = fifo_small_mix_cols_6_in_state_full;

assign fifo_small_mix_cols_7_in_state_data = shift_rows_8_out_state_data;
assign fifo_small_mix_cols_7_in_state_wr = shift_rows_8_out_state_wr;
assign shift_rows_8_out_state_full = fifo_small_mix_cols_7_in_state_full;

assign fifo_small_mix_cols_8_in_state_data = shift_rows_9_out_state_data;
assign fifo_small_mix_cols_8_in_state_wr = shift_rows_9_out_state_wr;
assign shift_rows_9_out_state_full = fifo_small_mix_cols_8_in_state_full;

endmodule
